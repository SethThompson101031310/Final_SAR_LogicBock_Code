// Created by ihdl
module SAR_FINAL_3(Q, array_gnd, array_vdd, comp_reg, data_clk_out, comp, compP, clk, rst_n,sh_clk, CAL_ext, CAL_out, PR_bar);


output [29:0] Q;
output array_gnd, array_vdd, data_clk_out, comp_reg, CAL_out, PR_bar;
input  comp, compP, clk, rst_n, sh_clk, CAL_ext;

// 'Cases'
parameter [4:0] INIT   = 5'b00000,
				CHARGE = 5'b00001,
                State9  = 5'b00011,
                State8  = 5'b00010,
                State7  = 5'b00110,
                State6  = 5'b00111,
                State5  = 5'b00101,
                State4  = 5'b00100,
                State3  = 5'b01100,
                State2  = 5'b01101,
                State1  = 5'b01111,
                State0  = 5'b01110,
                CAL1    = 5'b01010,
                CAL2    = 5'b01011,
                CAL3    = 5'b01001,
                CAL4    = 5'b01000,
                CAL5    = 5'b11000,
                RESET   = 5'b11001;

// 'States'
parameter [9:0] NONE     = 10'b0000000000,
                State9_1 = 10'b0000000001,
                State8_1 = 10'b0000000010,
                State8_3 = 10'b0000000011,
                State7_1 = 10'b0000000100,
                State7_3 = 10'b0000000101,
                State7_5 = 10'b0000000110,
                State7_7 = 10'b0000000111,
                State6_1 = 10'b0000001000,
                State6_3 = 10'b0000001001,
                State6_5 = 10'b0000001010,
                State6_7 = 10'b0000001011,
                State6_9 = 10'b0000001100,
                State6_11= 10'b0000001101,
                State6_13= 10'b0000001110,
                State6_15= 10'b0000001111,
                State5_1 = 10'b0000010000,
                State5_3 = 10'b0000010001,
                State5_5 = 10'b0000010010,
                State5_7 = 10'b0000010011,
                State5_9 = 10'b0000010100,
                State5_11= 10'b0000010101,
                State5_13= 10'b0000010110,
                State5_15= 10'b0000010111,
                State5_17= 10'b0000011000,
                State5_19= 10'b0000011001,
                State5_21= 10'b0000011010,
                State5_23= 10'b0000011011,
                State5_25= 10'b0000011100,
                State5_27= 10'b0000011101,
                State5_29= 10'b0000011110,
                State5_31= 10'b0000011111,
                State4_1 = 10'b0000100000,
                State4_3 = 10'b0000100001,
                State4_5 = 10'b0000100010,
                State4_7 = 10'b0000100011,
                State4_9 = 10'b0000100100,
                State4_11= 10'b0000100101,
                State4_13= 10'b0000100110,
                State4_15= 10'b0000100111,
                State4_17= 10'b0000101000,
                State4_19= 10'b0000101001,
                State4_21= 10'b0000101010,
                State4_23= 10'b0000101011,
                State4_25= 10'b0000101100,
                State4_27= 10'b0000101101,
                State4_29= 10'b0000101110,
                State4_31= 10'b0000101111,
                State4_33= 10'b0000110000,
                State4_35= 10'b0000110001,
                State4_37= 10'b0000110010,
                State4_39= 10'b0000110011,
                State4_41= 10'b0000110100,
                State4_43= 10'b0000110101,
                State4_45= 10'b0000110110,
                State4_47= 10'b0000110111,
                State4_49= 10'b0000111000,
                State4_51= 10'b0000111001,
                State4_53= 10'b0000111010,
                State4_55= 10'b0000111011,
                State4_57= 10'b0000111100,
                State4_59= 10'b0000111101,
                State4_61= 10'b0000111110,
                State4_63= 10'b0000111111,
                State3_1 = 10'b0001000000,
                State3_3 = 10'b0001000001,
                State3_5 = 10'b0001000010,
                State3_7 = 10'b0001000011,
                State3_9 = 10'b0001000100,
                State3_11= 10'b0001000101,
                State3_13= 10'b0001000110,
                State3_15= 10'b0001000111,
                State3_17= 10'b0001001000,
                State3_19= 10'b0001001001,
                State3_21= 10'b0001001010,
                State3_23= 10'b0001001011,
                State3_25= 10'b0001001100,
                State3_27= 10'b0001001101,
                State3_29= 10'b0001001110,
                State3_31= 10'b0001001111,
                State3_33= 10'b0001010000,
                State3_35= 10'b0001010001,
                State3_37= 10'b0001010010,
                State3_39= 10'b0001010011,
                State3_41= 10'b0001010100,
                State3_43= 10'b0001010101,
                State3_45= 10'b0001010110,
                State3_47= 10'b0001010111,
                State3_49= 10'b0001011000,
                State3_51= 10'b0001011001,
                State3_53= 10'b0001011010,
                State3_55= 10'b0001011011,
                State3_57= 10'b0001011100,
                State3_59= 10'b0001011101,
                State3_61= 10'b0001011110,
                State3_63= 10'b0001011111,
                State3_65= 10'b0001100000,
                State3_67= 10'b0001100001,
                State3_69= 10'b0001100010,
                State3_71= 10'b0001100011,
                State3_73= 10'b0001100100,
                State3_75= 10'b0001100101,
                State3_77= 10'b0001100110,
                State3_79= 10'b0001100111,
                State3_81= 10'b0001101000,
                State3_83= 10'b0001101001,
                State3_85= 10'b0001101010,
                State3_87= 10'b0001101011,
                State3_89= 10'b0001101100,
                State3_91= 10'b0001101101,
                State3_93= 10'b0001101110,
                State3_95= 10'b0001101111,
                State3_97= 10'b0001110000,
                State3_99= 10'b0001110001,
                State3_101= 10'b0001110010,
                State3_103= 10'b0001110011,
                State3_105= 10'b0001110100,
                State3_107= 10'b0001110101,
                State3_109= 10'b0001110110,
                State3_111= 10'b0001110111,
                State3_113= 10'b0001111000,
                State3_115= 10'b0001111001,
                State3_117= 10'b0001111010,
                State3_119= 10'b0001111011,
                State3_121= 10'b0001111100,
                State3_123= 10'b0001111101,
                State3_125= 10'b0001111110,
                State3_127= 10'b0001111111,
                State2_1 = 10'b0010000000,
                State2_3 = 10'b0010000001,
                State2_5 = 10'b0010000010,
                State2_7 = 10'b0010000011,
                State2_9 = 10'b0010000100,
                State2_11= 10'b0010000101,
                State2_13= 10'b0010000110,
                State2_15= 10'b0010000111,
                State2_17= 10'b0010001000,
                State2_19= 10'b0010001001,
                State2_21= 10'b0010001010,
                State2_23= 10'b0010001011,
                State2_25= 10'b0010001100,
                State2_27= 10'b0010001101,
                State2_29= 10'b0010001110,
                State2_31= 10'b0010001111,
                State2_33= 10'b0010010000,
                State2_35= 10'b0010010001,
                State2_37= 10'b0010010010,
                State2_39= 10'b0010010011,
                State2_41= 10'b0010010100,
                State2_43= 10'b0010010101,
                State2_45= 10'b0010010110,
                State2_47= 10'b0010010111,
                State2_49= 10'b0010011000,
                State2_51= 10'b0010011001,
                State2_53= 10'b0010011010,
                State2_55= 10'b0010011011,
                State2_57= 10'b0010011100,
                State2_59= 10'b0010011101,
                State2_61= 10'b0010011110,
                State2_63= 10'b0010011111,
                State2_65= 10'b0010100000,
                State2_67= 10'b0010100001,
                State2_69= 10'b0010100010,
                State2_71= 10'b0010100011,
                State2_73= 10'b0010100100,
                State2_75= 10'b0010100101,
                State2_77= 10'b0010100110,
                State2_79= 10'b0010100111,
                State2_81= 10'b0010101000,
                State2_83= 10'b0010101001,
                State2_85= 10'b0010101010,
                State2_87= 10'b0010101011,
                State2_89= 10'b0010101100,
                State2_91= 10'b0010101101,
                State2_93= 10'b0010101110,
                State2_95= 10'b0010101111,
                State2_97= 10'b0010110000,
                State2_99= 10'b0010110001,
                State2_101= 10'b0010110010,
                State2_103= 10'b0010110011,
                State2_105= 10'b0010110100,
                State2_107= 10'b0010110101,
                State2_109= 10'b0010110110,
                State2_111= 10'b0010110111,
                State2_113= 10'b0010111000,
                State2_115= 10'b0010111001,
                State2_117= 10'b0010111010,
                State2_119= 10'b0010111011,
                State2_121= 10'b0010111100,
                State2_123= 10'b0010111101,
                State2_125= 10'b0010111110,
                State2_127= 10'b0010111111,
                State2_129= 10'b0011000000,
                State2_131= 10'b0011000001,
                State2_133= 10'b0011000010,
                State2_135= 10'b0011000011,
                State2_137= 10'b0011000100,
                State2_139= 10'b0011000101,
                State2_141= 10'b0011000110,
                State2_143= 10'b0011000111,
                State2_145= 10'b0011001000,
                State2_147= 10'b0011001001,
                State2_149= 10'b0011001010,
                State2_151= 10'b0011001011,
                State2_153= 10'b0011001100,
                State2_155= 10'b0011001101,
                State2_157= 10'b0011001110,
                State2_159= 10'b0011001111,
                State2_161= 10'b0011010000,
                State2_163= 10'b0011010001,
                State2_165= 10'b0011010010,
                State2_167= 10'b0011010011,
                State2_169= 10'b0011010100,
                State2_171= 10'b0011010101,
                State2_173= 10'b0011010110,
                State2_175= 10'b0011010111,
                State2_177= 10'b0011011000,
                State2_179= 10'b0011011001,
                State2_181= 10'b0011011010,
                State2_183= 10'b0011011011,
                State2_185= 10'b0011011100,
                State2_187= 10'b0011011101,
                State2_189= 10'b0011011110,
                State2_191= 10'b0011011111,
                State2_193= 10'b0011100000,
                State2_195= 10'b0011100001,
                State2_197= 10'b0011100010,
                State2_199= 10'b0011100011,
                State2_201= 10'b0011100100,
                State2_203= 10'b0011100101,
                State2_205= 10'b0011100110,
                State2_207= 10'b0011100111,
                State2_209= 10'b0011101000,
                State2_211= 10'b0011101001,
                State2_213= 10'b0011101010,
                State2_215= 10'b0011101011,
                State2_217= 10'b0011101100,
                State2_219= 10'b0011101101,
                State2_221= 10'b0011101110,
                State2_223= 10'b0011101111,
                State2_225= 10'b0011110000,
                State2_227= 10'b0011110001,
                State2_229= 10'b0011110010,
                State2_231= 10'b0011110011,
                State2_233= 10'b0011110100,
                State2_235= 10'b0011110101,
                State2_237= 10'b0011110110,
                State2_239= 10'b0011110111,
                State2_241= 10'b0011111000,
                State2_243= 10'b0011111001,
                State2_245= 10'b0011111010,
                State2_247= 10'b0011111011,
                State2_249= 10'b0011111100,
                State2_251= 10'b0011111101,
                State2_253= 10'b0011111110,
                State2_255= 10'b0011111111,
                State1_1 = 10'b0100000000,
                State1_3 = 10'b0100000001,
                State1_5 = 10'b0100000010,
                State1_7 = 10'b0100000011,
                State1_9 = 10'b0100000100,
                State1_11= 10'b0100000101,
                State1_13= 10'b0100000110,
                State1_15= 10'b0100000111,
                State1_17= 10'b0100001000,
                State1_19= 10'b0100001001,
                State1_21= 10'b0100001010,
                State1_23= 10'b0100001011,
                State1_25= 10'b0100001100,
                State1_27= 10'b0100001101,
                State1_29= 10'b0100001110,
                State1_31= 10'b0100001111,
                State1_33= 10'b0100010000,
                State1_35= 10'b0100010001,
                State1_37= 10'b0100010010,
                State1_39= 10'b0100010011,
                State1_41= 10'b0100010100,
                State1_43= 10'b0100010101,
                State1_45= 10'b0100010110,
                State1_47= 10'b0100010111,
                State1_49= 10'b0100011000,
                State1_51= 10'b0100011001,
                State1_53= 10'b0100011010,
                State1_55= 10'b0100011011,
                State1_57= 10'b0100011100,
                State1_59= 10'b0100011101,
                State1_61= 10'b0100011110,
                State1_63= 10'b0100011111,
                State1_65= 10'b0100100000,
                State1_67= 10'b0100100001,
                State1_69= 10'b0100100010,
                State1_71= 10'b0100100011,
                State1_73= 10'b0100100100,
                State1_75= 10'b0100100101,
                State1_77= 10'b0100100110,
                State1_79= 10'b0100100111,
                State1_81= 10'b0100101000,
                State1_83= 10'b0100101001,
                State1_85= 10'b0100101010,
                State1_87= 10'b0100101011,
                State1_89= 10'b0100101100,
                State1_91= 10'b0100101101,
                State1_93= 10'b0100101110,
                State1_95= 10'b0100101111,
                State1_97= 10'b0100110000,
                State1_99= 10'b0100110001,
                State1_101= 10'b0100110010,
                State1_103= 10'b0100110011,
                State1_105= 10'b0100110100,
                State1_107= 10'b0100110101,
                State1_109= 10'b0100110110,
                State1_111= 10'b0100110111,
                State1_113= 10'b0100111000,
                State1_115= 10'b0100111001,
                State1_117= 10'b0100111010,
                State1_119= 10'b0100111011,
                State1_121= 10'b0100111100,
                State1_123= 10'b0100111101,
                State1_125= 10'b0100111110,
                State1_127= 10'b0100111111,
                State1_129= 10'b0101000000,
                State1_131= 10'b0101000001,
                State1_133= 10'b0101000010,
                State1_135= 10'b0101000011,
                State1_137= 10'b0101000100,
                State1_139= 10'b0101000101,
                State1_141= 10'b0101000110,
                State1_143= 10'b0101000111,
                State1_145= 10'b0101001000,
                State1_147= 10'b0101001001,
                State1_149= 10'b0101001010,
                State1_151= 10'b0101001011,
                State1_153= 10'b0101001100,
                State1_155= 10'b0101001101,
                State1_157= 10'b0101001110,
                State1_159= 10'b0101001111,
                State1_161= 10'b0101010000,
                State1_163= 10'b0101010001,
                State1_165= 10'b0101010010,
                State1_167= 10'b0101010011,
                State1_169= 10'b0101010100,
                State1_171= 10'b0101010101,
                State1_173= 10'b0101010110,
                State1_175= 10'b0101010111,
                State1_177= 10'b0101011000,
                State1_179= 10'b0101011001,
                State1_181= 10'b0101011010,
                State1_183= 10'b0101011011,
                State1_185= 10'b0101011100,
                State1_187= 10'b0101011101,
                State1_189= 10'b0101011110,
                State1_191= 10'b0101011111,
                State1_193= 10'b0101100000,
                State1_195= 10'b0101100001,
                State1_197= 10'b0101100010,
                State1_199= 10'b0101100011,
                State1_201= 10'b0101100100,
                State1_203= 10'b0101100101,
                State1_205= 10'b0101100110,
                State1_207= 10'b0101100111,
                State1_209= 10'b0101101000,
                State1_211= 10'b0101101001,
                State1_213= 10'b0101101010,
                State1_215= 10'b0101101011,
                State1_217= 10'b0101101100,
                State1_219= 10'b0101101101,
                State1_221= 10'b0101101110,
                State1_223= 10'b0101101111,
                State1_225= 10'b0101110000,
                State1_227= 10'b0101110001,
                State1_229= 10'b0101110010,
                State1_231= 10'b0101110011,
                State1_233= 10'b0101110100,
                State1_235= 10'b0101110101,
                State1_237= 10'b0101110110,
                State1_239= 10'b0101110111,
                State1_241= 10'b0101111000,
                State1_243= 10'b0101111001,
                State1_245= 10'b0101111010,
                State1_247= 10'b0101111011,
                State1_249= 10'b0101111100,
                State1_251= 10'b0101111101,
                State1_253= 10'b0101111110,
                State1_255= 10'b0101111111,
                State1_257= 10'b0110000000,
                State1_259= 10'b0110000001,
                State1_261= 10'b0110000010,
                State1_263= 10'b0110000011,
                State1_265= 10'b0110000100,
                State1_267= 10'b0110000101,
                State1_269= 10'b0110000110,
                State1_271= 10'b0110000111,
                State1_273= 10'b0110001000,
                State1_275= 10'b0110001001,
                State1_277= 10'b0110001010,
                State1_279= 10'b0110001011,
                State1_281= 10'b0110001100,
                State1_283= 10'b0110001101,
                State1_285= 10'b0110001110,
                State1_287= 10'b0110001111,
                State1_289= 10'b0110010000,
                State1_291= 10'b0110010001,
                State1_293= 10'b0110010010,
                State1_295= 10'b0110010011,
                State1_297= 10'b0110010100,
                State1_299= 10'b0110010101,
                State1_301= 10'b0110010110,
                State1_303= 10'b0110010111,
                State1_305= 10'b0110011000,
                State1_307= 10'b0110011001,
                State1_309= 10'b0110011010,
                State1_311= 10'b0110011011,
                State1_313= 10'b0110011100,
                State1_315= 10'b0110011101,
                State1_317= 10'b0110011110,
                State1_319= 10'b0110011111,
                State1_321= 10'b0110100000,
                State1_323= 10'b0110100001,
                State1_325= 10'b0110100010,
                State1_327= 10'b0110100011,
                State1_329= 10'b0110100100,
                State1_331= 10'b0110100101,
                State1_333= 10'b0110100110,
                State1_335= 10'b0110100111,
                State1_337= 10'b0110101000,
                State1_339= 10'b0110101001,
                State1_341= 10'b0110101010,
                State1_343= 10'b0110101011,
                State1_345= 10'b0110101100,
                State1_347= 10'b0110101101,
                State1_349= 10'b0110101110,
                State1_351= 10'b0110101111,
                State1_353= 10'b0110110000,
                State1_355= 10'b0110110001,
                State1_357= 10'b0110110010,
                State1_359= 10'b0110110011,
                State1_361= 10'b0110110100,
                State1_363= 10'b0110110101,
                State1_365= 10'b0110110110,
                State1_367= 10'b0110110111,
                State1_369= 10'b0110111000,
                State1_371= 10'b0110111001,
                State1_373= 10'b0110111010,
                State1_375= 10'b0110111011,
                State1_377= 10'b0110111100,
                State1_379= 10'b0110111101,
                State1_381= 10'b0110111110,
                State1_383= 10'b0110111111,
                State1_385= 10'b0111000000,
                State1_387= 10'b0111000001,
                State1_389= 10'b0111000010,
                State1_391= 10'b0111000011,
                State1_393= 10'b0111000100,
                State1_395= 10'b0111000101,
                State1_397= 10'b0111000110,
                State1_399= 10'b0111000111,
                State1_401= 10'b0111001000,
                State1_403= 10'b0111001001,
                State1_405= 10'b0111001010,
                State1_407= 10'b0111001011,
                State1_409= 10'b0111001100,
                State1_411= 10'b0111001101,
                State1_413= 10'b0111001110,
                State1_415= 10'b0111001111,
                State1_417= 10'b0111010000,
                State1_419= 10'b0111010001,
                State1_421= 10'b0111010010,
                State1_423= 10'b0111010011,
                State1_425= 10'b0111010100,
                State1_427= 10'b0111010101,
                State1_429= 10'b0111010110,
                State1_431= 10'b0111010111,
                State1_433= 10'b0111011000,
                State1_435= 10'b0111011001,
                State1_437= 10'b0111011010,
                State1_439= 10'b0111011011,
                State1_441= 10'b0111011100,
                State1_443= 10'b0111011101,
                State1_445= 10'b0111011110,
                State1_447= 10'b0111011111,
                State1_449= 10'b0111100000,
                State1_451= 10'b0111100001,
                State1_453= 10'b0111100010,
                State1_455= 10'b0111100011,
                State1_457= 10'b0111100100,
                State1_459= 10'b0111100101,
                State1_461= 10'b0111100110,
                State1_463= 10'b0111100111,
                State1_465= 10'b0111101000,
                State1_467= 10'b0111101001,
                State1_469= 10'b0111101010,
                State1_471= 10'b0111101011,
                State1_473= 10'b0111101100,
                State1_475= 10'b0111101101,
                State1_477= 10'b0111101110,
                State1_479= 10'b0111101111,
                State1_481= 10'b0111110000,
                State1_483= 10'b0111110001,
                State1_485= 10'b0111110010,
                State1_487= 10'b0111110011,
                State1_489= 10'b0111110100,
                State1_491= 10'b0111110101,
                State1_493= 10'b0111110110,
                State1_495= 10'b0111110111,
                State1_497= 10'b0111111000,
                State1_499= 10'b0111111001,
                State1_501= 10'b0111111010,
                State1_503= 10'b0111111011,
                State1_505= 10'b0111111100,
                State1_507= 10'b0111111101,
                State1_509= 10'b0111111110,
                State1_511= 10'b0111111111,
                State0_1 = 10'b1000000000,
                State0_3 = 10'b1000000001,
                State0_5 = 10'b1000000010,
                State0_7 = 10'b1000000011,
                State0_9 = 10'b1000000100,
                State0_11= 10'b1000000101,
                State0_13= 10'b1000000110,
                State0_15= 10'b1000000111,
                State0_17= 10'b1000001000,
                State0_19= 10'b1000001001,
                State0_21= 10'b1000001010,
                State0_23= 10'b1000001011,
                State0_25= 10'b1000001100,
                State0_27= 10'b1000001101,
                State0_29= 10'b1000001110,
                State0_31= 10'b1000001111,
                State0_33= 10'b1000010000,
                State0_35= 10'b1000010001,
                State0_37= 10'b1000010010,
                State0_39= 10'b1000010011,
                State0_41= 10'b1000010100,
                State0_43= 10'b1000010101,
                State0_45= 10'b1000010110,
                State0_47= 10'b1000010111,
                State0_49= 10'b1000011000,
                State0_51= 10'b1000011001,
                State0_53= 10'b1000011010,
                State0_55= 10'b1000011011,
                State0_57= 10'b1000011100,
                State0_59= 10'b1000011101,
                State0_61= 10'b1000011110,
                State0_63= 10'b1000011111,
                State0_65= 10'b1000100000,
                State0_67= 10'b1000100001,
                State0_69= 10'b1000100010,
                State0_71= 10'b1000100011,
                State0_73= 10'b1000100100,
                State0_75= 10'b1000100101,
                State0_77= 10'b1000100110,
                State0_79= 10'b1000100111,
                State0_81= 10'b1000101000,
                State0_83= 10'b1000101001,
                State0_85= 10'b1000101010,
                State0_87= 10'b1000101011,
                State0_89= 10'b1000101100,
                State0_91= 10'b1000101101,
                State0_93= 10'b1000101110,
                State0_95= 10'b1000101111,
                State0_97= 10'b1000110000,
                State0_99= 10'b1000110001,
                State0_101= 10'b1000110010,
                State0_103= 10'b1000110011,
                State0_105= 10'b1000110100,
                State0_107= 10'b1000110101,
                State0_109= 10'b1000110110,
                State0_111= 10'b1000110111,
                State0_113= 10'b1000111000,
                State0_115= 10'b1000111001,
                State0_117= 10'b1000111010,
                State0_119= 10'b1000111011,
                State0_121= 10'b1000111100,
                State0_123= 10'b1000111101,
                State0_125= 10'b1000111110,
                State0_127= 10'b1000111111,
                State0_129= 10'b1001000000,
                State0_131= 10'b1001000001,
                State0_133= 10'b1001000010,
                State0_135= 10'b1001000011,
                State0_137= 10'b1001000100,
                State0_139= 10'b1001000101,
                State0_141= 10'b1001000110,
                State0_143= 10'b1001000111,
                State0_145= 10'b1001001000,
                State0_147= 10'b1001001001,
                State0_149= 10'b1001001010,
                State0_151= 10'b1001001011,
                State0_153= 10'b1001001100,
                State0_155= 10'b1001001101,
                State0_157= 10'b1001001110,
                State0_159= 10'b1001001111,
                State0_161= 10'b1001010000,
                State0_163= 10'b1001010001,
                State0_165= 10'b1001010010,
                State0_167= 10'b1001010011,
                State0_169= 10'b1001010100,
                State0_171= 10'b1001010101,
                State0_173= 10'b1001010110,
                State0_175= 10'b1001010111,
                State0_177= 10'b1001011000,
                State0_179= 10'b1001011001,
                State0_181= 10'b1001011010,
                State0_183= 10'b1001011011,
                State0_185= 10'b1001011100,
                State0_187= 10'b1001011101,
                State0_189= 10'b1001011110,
                State0_191= 10'b1001011111,
                State0_193= 10'b1001100000,
                State0_195= 10'b1001100001,
                State0_197= 10'b1001100010,
                State0_199= 10'b1001100011,
                State0_201= 10'b1001100100,
                State0_203= 10'b1001100101,
                State0_205= 10'b1001100110,
                State0_207= 10'b1001100111,
                State0_209= 10'b1001101000,
                State0_211= 10'b1001101001,
                State0_213= 10'b1001101010,
                State0_215= 10'b1001101011,
                State0_217= 10'b1001101100,
                State0_219= 10'b1001101101,
                State0_221= 10'b1001101110,
                State0_223= 10'b1001101111,
                State0_225= 10'b1001110000,
                State0_227= 10'b1001110001,
                State0_229= 10'b1001110010,
                State0_231= 10'b1001110011,
                State0_233= 10'b1001110100,
                State0_235= 10'b1001110101,
                State0_237= 10'b1001110110,
                State0_239= 10'b1001110111,
                State0_241= 10'b1001111000,
                State0_243= 10'b1001111001,
                State0_245= 10'b1001111010,
                State0_247= 10'b1001111011,
                State0_249= 10'b1001111100,
                State0_251= 10'b1001111101,
                State0_253= 10'b1001111110,
                State0_255= 10'b1001111111,
                State0_257= 10'b1010000000,
                State0_259= 10'b1010000001,
                State0_261= 10'b1010000010,
                State0_263= 10'b1010000011,
                State0_265= 10'b1010000100,
                State0_267= 10'b1010000101,
                State0_269= 10'b1010000110,
                State0_271= 10'b1010000111,
                State0_273= 10'b1010001000,
                State0_275= 10'b1010001001,
                State0_277= 10'b1010001010,
                State0_279= 10'b1010001011,
                State0_281= 10'b1010001100,
                State0_283= 10'b1010001101,
                State0_285= 10'b1010001110,
                State0_287= 10'b1010001111,
                State0_289= 10'b1010010000,
                State0_291= 10'b1010010001,
                State0_293= 10'b1010010010,
                State0_295= 10'b1010010011,
                State0_297= 10'b1010010100,
                State0_299= 10'b1010010101,
                State0_301= 10'b1010010110,
                State0_303= 10'b1010010111,
                State0_305= 10'b1010011000,
                State0_307= 10'b1010011001,
                State0_309= 10'b1010011010,
                State0_311= 10'b1010011011,
                State0_313= 10'b1010011100,
                State0_315= 10'b1010011101,
                State0_317= 10'b1010011110,
                State0_319= 10'b1010011111,
                State0_321= 10'b1010100000,
                State0_323= 10'b1010100001,
                State0_325= 10'b1010100010,
                State0_327= 10'b1010100011,
                State0_329= 10'b1010100100,
                State0_331= 10'b1010100101,
                State0_333= 10'b1010100110,
                State0_335= 10'b1010100111,
                State0_337= 10'b1010101000,
                State0_339= 10'b1010101001,
                State0_341= 10'b1010101010,
                State0_343= 10'b1010101011,
                State0_345= 10'b1010101100,
                State0_347= 10'b1010101101,
                State0_349= 10'b1010101110,
                State0_351= 10'b1010101111,
                State0_353= 10'b1010110000,
                State0_355= 10'b1010110001,
                State0_357= 10'b1010110010,
                State0_359= 10'b1010110011,
                State0_361= 10'b1010110100,
                State0_363= 10'b1010110101,
                State0_365= 10'b1010110110,
                State0_367= 10'b1010110111,
                State0_369= 10'b1010111000,
                State0_371= 10'b1010111001,
                State0_373= 10'b1010111010,
                State0_375= 10'b1010111011,
                State0_377= 10'b1010111100,
                State0_379= 10'b1010111101,
                State0_381= 10'b1010111110,
                State0_383= 10'b1010111111,
                State0_385= 10'b1011000000,
                State0_387= 10'b1011000001,
                State0_389= 10'b1011000010,
                State0_391= 10'b1011000011,
                State0_393= 10'b1011000100,
                State0_395= 10'b1011000101,
                State0_397= 10'b1011000110,
                State0_399= 10'b1011000111,
                State0_401= 10'b1011001000,
                State0_403= 10'b1011001001,
                State0_405= 10'b1011001010,
                State0_407= 10'b1011001011,
                State0_409= 10'b1011001100,
                State0_411= 10'b1011001101,
                State0_413= 10'b1011001110,
                State0_415= 10'b1011001111,
                State0_417= 10'b1011010000,
                State0_419= 10'b1011010001,
                State0_421= 10'b1011010010,
                State0_423= 10'b1011010011,
                State0_425= 10'b1011010100,
                State0_427= 10'b1011010101,
                State0_429= 10'b1011010110,
                State0_431= 10'b1011010111,
                State0_433= 10'b1011011000,
                State0_435= 10'b1011011001,
                State0_437= 10'b1011011010,
                State0_439= 10'b1011011011,
                State0_441= 10'b1011011100,
                State0_443= 10'b1011011101,
                State0_445= 10'b1011011110,
                State0_447= 10'b1011011111,
                State0_449= 10'b1011100000,
                State0_451= 10'b1011100001,
                State0_453= 10'b1011100010,
                State0_455= 10'b1011100011,
                State0_457= 10'b1011100100,
                State0_459= 10'b1011100101,
                State0_461= 10'b1011100110,
                State0_463= 10'b1011100111,
                State0_465= 10'b1011101000,
                State0_467= 10'b1011101001,
                State0_469= 10'b1011101010,
                State0_471= 10'b1011101011,
                State0_473= 10'b1011101100,
                State0_475= 10'b1011101101,
                State0_477= 10'b1011101110,
                State0_479= 10'b1011101111,
                State0_481= 10'b1011110000,
                State0_483= 10'b1011110001,
                State0_485= 10'b1011110010,
                State0_487= 10'b1011110011,
                State0_489= 10'b1011110100,
                State0_491= 10'b1011110101,
                State0_493= 10'b1011110110,
                State0_495= 10'b1011110111,
                State0_497= 10'b1011111000,
                State0_499= 10'b1011111001,
                State0_501= 10'b1011111010,
                State0_503= 10'b1011111011,
                State0_505= 10'b1011111100,
                State0_507= 10'b1011111101,
                State0_509= 10'b1011111110,
                State0_511= 10'b1011111111,
                State0_513= 10'b1100000000,
                State0_515= 10'b1100000001,
                State0_517= 10'b1100000010,
                State0_519= 10'b1100000011,
                State0_521= 10'b1100000100,
                State0_523= 10'b1100000101,
                State0_525= 10'b1100000110,
                State0_527= 10'b1100000111,
                State0_529= 10'b1100001000,
                State0_531= 10'b1100001001,
                State0_533= 10'b1100001010,
                State0_535= 10'b1100001011,
                State0_537= 10'b1100001100,
                State0_539= 10'b1100001101,
                State0_541= 10'b1100001110,
                State0_543= 10'b1100001111,
                State0_545= 10'b1100010000,
                State0_547= 10'b1100010001,
                State0_549= 10'b1100010010,
                State0_551= 10'b1100010011,
                State0_553= 10'b1100010100,
                State0_555= 10'b1100010101,
                State0_557= 10'b1100010110,
                State0_559= 10'b1100010111,
                State0_561= 10'b1100011000,
                State0_563= 10'b1100011001,
                State0_565= 10'b1100011010,
                State0_567= 10'b1100011011,
                State0_569= 10'b1100011100,
                State0_571= 10'b1100011101,
                State0_573= 10'b1100011110,
                State0_575= 10'b1100011111,
                State0_577= 10'b1100100000,
                State0_579= 10'b1100100001,
                State0_581= 10'b1100100010,
                State0_583= 10'b1100100011,
                State0_585= 10'b1100100100,
                State0_587= 10'b1100100101,
                State0_589= 10'b1100100110,
                State0_591= 10'b1100100111,
                State0_593= 10'b1100101000,
                State0_595= 10'b1100101001,
                State0_597= 10'b1100101010,
                State0_599= 10'b1100101011,
                State0_601= 10'b1100101100,
                State0_603= 10'b1100101101,
                State0_605= 10'b1100101110,
                State0_607= 10'b1100101111,
                State0_609= 10'b1100110000,
                State0_611= 10'b1100110001,
                State0_613= 10'b1100110010,
                State0_615= 10'b1100110011,
                State0_617= 10'b1100110100,
                State0_619= 10'b1100110101,
                State0_621= 10'b1100110110,
                State0_623= 10'b1100110111,
                State0_625= 10'b1100111000,
                State0_627= 10'b1100111001,
                State0_629= 10'b1100111010,
                State0_631= 10'b1100111011,
                State0_633= 10'b1100111100,
                State0_635= 10'b1100111101,
                State0_637= 10'b1100111110,
                State0_639= 10'b1100111111,
                State0_641= 10'b1101000000,
                State0_643= 10'b1101000001,
                State0_645= 10'b1101000010,
                State0_647= 10'b1101000011,
                State0_649= 10'b1101000100,
                State0_651= 10'b1101000101,
                State0_653= 10'b1101000110,
                State0_655= 10'b1101000111,
                State0_657= 10'b1101001000,
                State0_659= 10'b1101001001,
                State0_661= 10'b1101001010,
                State0_663= 10'b1101001011,
                State0_665= 10'b1101001100,
                State0_667= 10'b1101001101,
                State0_669= 10'b1101001110,
                State0_671= 10'b1101001111,
                State0_673= 10'b1101010000,
                State0_675= 10'b1101010001,
                State0_677= 10'b1101010010,
                State0_679= 10'b1101010011,
                State0_681= 10'b1101010100,
                State0_683= 10'b1101010101,
                State0_685= 10'b1101010110,
                State0_687= 10'b1101010111,
                State0_689= 10'b1101011000,
                State0_691= 10'b1101011001,
                State0_693= 10'b1101011010,
                State0_695= 10'b1101011011,
                State0_697= 10'b1101011100,
                State0_699= 10'b1101011101,
                State0_701= 10'b1101011110,
                State0_703= 10'b1101011111,
                State0_705= 10'b1101100000,
                State0_707= 10'b1101100001,
                State0_709= 10'b1101100010,
                State0_711= 10'b1101100011,
                State0_713= 10'b1101100100,
                State0_715= 10'b1101100101,
                State0_717= 10'b1101100110,
                State0_719= 10'b1101100111,
                State0_721= 10'b1101101000,
                State0_723= 10'b1101101001,
                State0_725= 10'b1101101010,
                State0_727= 10'b1101101011,
                State0_729= 10'b1101101100,
                State0_731= 10'b1101101101,
                State0_733= 10'b1101101110,
                State0_735= 10'b1101101111,
                State0_737= 10'b1101110000,
                State0_739= 10'b1101110001,
                State0_741= 10'b1101110010,
                State0_743= 10'b1101110011,
                State0_745= 10'b1101110100,
                State0_747= 10'b1101110101,
                State0_749= 10'b1101110110,
                State0_751= 10'b1101110111,
                State0_753= 10'b1101111000,
                State0_755= 10'b1101111001,
                State0_757= 10'b1101111010,
                State0_759= 10'b1101111011,
                State0_761= 10'b1101111100,
                State0_763= 10'b1101111101,
                State0_765= 10'b1101111110,
                State0_767= 10'b1101111111,
                State0_769= 10'b1110000000,
                State0_771= 10'b1110000001,
                State0_773= 10'b1110000010,
                State0_775= 10'b1110000011,
                State0_777= 10'b1110000100,
                State0_779= 10'b1110000101,
                State0_781= 10'b1110000110,
                State0_783= 10'b1110000111,
                State0_785= 10'b1110001000,
                State0_787= 10'b1110001001,
                State0_789= 10'b1110001010,
                State0_791= 10'b1110001011,
                State0_793= 10'b1110001100,
                State0_795= 10'b1110001101,
                State0_797= 10'b1110001110,
                State0_799= 10'b1110001111,
                State0_801= 10'b1110010000,
                State0_803= 10'b1110010001,
                State0_805= 10'b1110010010,
                State0_807= 10'b1110010011,
                State0_809= 10'b1110010100,
                State0_811= 10'b1110010101,
                State0_813= 10'b1110010110,
                State0_815= 10'b1110010111,
                State0_817= 10'b1110011000,
                State0_819= 10'b1110011001,
                State0_821= 10'b1110011010,
                State0_823= 10'b1110011011,
                State0_825= 10'b1110011100,
                State0_827= 10'b1110011101,
                State0_829= 10'b1110011110,
                State0_831= 10'b1110011111,
                State0_833= 10'b1110100000,
                State0_835= 10'b1110100001,
                State0_837= 10'b1110100010,
                State0_839= 10'b1110100011,
                State0_841= 10'b1110100100,
                State0_843= 10'b1110100101,
                State0_845= 10'b1110100110,
                State0_847= 10'b1110100111,
                State0_849= 10'b1110101000,
                State0_851= 10'b1110101001,
                State0_853= 10'b1110101010,
                State0_855= 10'b1110101011,
                State0_857= 10'b1110101100,
                State0_859= 10'b1110101101,
                State0_861= 10'b1110101110,
                State0_863= 10'b1110101111,
                State0_865= 10'b1110110000,
                State0_867= 10'b1110110001,
                State0_869= 10'b1110110010,
                State0_871= 10'b1110110011,
                State0_873= 10'b1110110100,
                State0_875= 10'b1110110101,
                State0_877= 10'b1110110110,
                State0_879= 10'b1110110111,
                State0_881= 10'b1110111000,
                State0_883= 10'b1110111001,
                State0_885= 10'b1110111010,
                State0_887= 10'b1110111011,
                State0_889= 10'b1110111100,
                State0_891= 10'b1110111101,
                State0_893= 10'b1110111110,
                State0_895= 10'b1110111111,
                State0_897= 10'b1111000000,
                State0_899= 10'b1111000001,
                State0_901= 10'b1111000010,
                State0_903= 10'b1111000011,
                State0_905= 10'b1111000100,
                State0_907= 10'b1111000101,
                State0_909= 10'b1111000110,
                State0_911= 10'b1111000111,
                State0_913= 10'b1111001000,
                State0_915= 10'b1111001001,
                State0_917= 10'b1111001010,
                State0_919= 10'b1111001011,
                State0_921= 10'b1111001100,
                State0_923= 10'b1111001101,
                State0_925= 10'b1111001110,
                State0_927= 10'b1111001111,
                State0_929= 10'b1111010000,
                State0_931= 10'b1111010001,
                State0_933= 10'b1111010010,
                State0_935= 10'b1111010011,
                State0_937= 10'b1111010100,
                State0_939= 10'b1111010101,
                State0_941= 10'b1111010110,
                State0_943= 10'b1111010111,
                State0_945= 10'b1111011000,
                State0_947= 10'b1111011001,
                State0_949= 10'b1111011010,
                State0_951= 10'b1111011011,
                State0_953= 10'b1111011100,
                State0_955= 10'b1111011101,
                State0_957= 10'b1111011110,
                State0_959= 10'b1111011111,
                State0_961= 10'b1111100000,
                State0_963= 10'b1111100001,
                State0_965= 10'b1111100010,
                State0_967= 10'b1111100011,
                State0_969= 10'b1111100100,
                State0_971= 10'b1111100101,
                State0_973= 10'b1111100110,
                State0_975= 10'b1111100111,
                State0_977= 10'b1111101000,
                State0_979= 10'b1111101001,
                State0_981= 10'b1111101010,
                State0_983= 10'b1111101011,
                State0_985= 10'b1111101100,
                State0_987= 10'b1111101101,
                State0_989= 10'b1111101110,
                State0_991= 10'b1111101111,
                State0_993= 10'b1111110000,
                State0_995= 10'b1111110001,
                State0_997= 10'b1111110010,
                State0_999= 10'b1111110011,
                State0_1001= 10'b1111110100,
                State0_1003= 10'b1111110101,
                State0_1005= 10'b1111110110,
                State0_1007= 10'b1111110111,
                State0_1009= 10'b1111111000,
                State0_1011= 10'b1111111001,
                State0_1013= 10'b1111111010,
                State0_1015= 10'b1111111011,
                State0_1017= 10'b1111111100,
                State0_1019= 10'b1111111101,
                State0_1021= 10'b1111111110,
                State0_1023= 10'b1111111111;

reg [4:0]   state;
reg [4:0]   next_state;
reg [9:0]   prev_state_reg;
reg [9:0]   prev_state;
reg [29:0]  Q;
reg [29:0]  Q_reg;
reg         array_vdd;
reg         array_gnd;
reg         data_clk_out;
reg         data_clk;
reg         comp_reg;
reg         get_comp;
reg         CAL_out;
reg         PR_bar;


always @ (negedge clk or negedge rst_n) begin
  if (!rst_n)
    begin
      state           <= RESET;
      prev_state_reg  <= NONE;
      comp_reg        <= 1'b0;
      data_clk_out    <= 1'b0;
    end
  else
    begin
      Q_reg  <= Q;
      if (sh_clk || CAL_ext)
         state          <= next_state;
      else
         state          <= INIT;
         prev_state_reg <= prev_state;
         data_clk_out   <= data_clk;

      if (get_comp)
         comp_reg       <= comp;
    end
end

always @ (state or comp or compP) begin

  if (clk && (!comp || !compP) && sh_clk) begin  
	Q = 30'b000000000000000000000000000000;
    array_vdd    = 1'b1;
    array_gnd    = 1'b0;
  end else begin

  // DEFAULT VALUES
  Q  = Q_reg;
  array_gnd     = 1'b0;
  array_vdd     = 1'b1;
  next_state    = INIT;
  prev_state    = prev_state_reg;
  data_clk      = 1'b0;
  get_comp      = 1'b0;
  PR_bar        = 1'b1;
  CAL_out       = 1'b0;

  case (state)
  RESET:
    begin
      next_state = INIT;
      Q = 30'b111111111111111111111111111111;
      array_gnd = 1'b1;
      array_vdd = 1'b1;
      CAL_out   = 1'b0;
      PR_bar    = 1'b1;
    end
  INIT:
    begin
      next_state = CHARGE;
      // When we initialize, first discharge all caps
	  // Only half need to be discharged since next state sets other half to 1
      Q = 30'b111111111111111000000000000000;
      array_gnd = 1'b1;
      array_vdd = 1'b1;
    end
  CHARGE:
    begin
	if (CAL_ext) begin
      next_state = CAL1;
      PR_bar     = 1'b0;
    end
    else
      next_state = State9;
      // Charge half the caps to 1
      Q = 30'b000000000000000111111111111111;
      array_gnd = 1'b0;
      array_vdd = 1'b0;
    end

// 5 STEP CALIBRATION
    CAL1:
      begin
        next_state = CAL2;
        Q = 30'b110000000000000110000000000000;
        CAL_out    = 1'b1;
        end
    CAL2:
      begin
        next_state = CAL3;
        Q = 30'b110000000000000110000000000000;
        CAL_out    = 1'b1;
        end
    CAL3:
      begin
        next_state = CAL4;
        Q = 30'b110000000000000110000000000000;
        CAL_out    = 1'b1;
        end
    CAL4:
      begin
        next_state = CAL5;
        Q = 30'b110000000000000110000000000000;
        CAL_out    = 1'b1;
        end
    CAL5:
      begin
        next_state = INIT;
        Q = 30'b110000000000000110000000000000;
        CAL_out    = 1'b1;
        end
  //////////////////
  
  State9:
    begin
		next_state = State8;
		data_clk = 1'b1;
        get_comp = 1'b1;
        // Must create 1/2*Vdd
        Q = 30'b110000000000000110000000000000;
	end
  State8:
    begin
        next_state = State7;
        data_clk = 1'b1;
        get_comp = 1'b1;
        if (comp_reg == 1'b0)
            begin
                // Must create 1/4*Vdd
                Q = 30'b111100000000000000000000000000;
                prev_state = State8_1;
            end
        if (comp_reg == 1'b1)
            begin
                // Must create 3/4*Vdd
                Q = 30'b110000000000000001100000000000;
                prev_state = State8_3;
            end
    end
  State7:
    begin
        next_state = State6;
        data_clk = 1'b1;
        get_comp = 1'b1;
        if (comp_reg == 1'b0 && prev_state_reg == State8_1)
            begin
                // Must create 1/8*Vdd
                Q = 30'b100010000000000000000000000000;
                prev_state = State7_1;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State8_1)
            begin
                // Must create 3/8*Vdd
                Q = 30'b100011100000000001100000000000;
                prev_state = State7_3;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State8_3)
            begin
                // Must create 5/8*Vdd
                Q = 30'b101100000000000000011100000000;
                prev_state = State7_5;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State8_3)
            begin
                // Must create 7/8*Vdd
                Q = 30'b100000000000000000010000000000;
                prev_state = State7_7;
            end
    end
  State6:
    begin
        next_state = State5;
        data_clk = 1'b1;
        get_comp = 1'b1;
        if (comp_reg == 1'b0 && prev_state_reg == State7_1)
            begin
                // Must create 1/16*Vdd
                Q = 30'b010001110000000000000000000000;
                prev_state = State6_1;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State7_1)
            begin
                // Must create 3/16*Vdd
                Q = 30'b100001111000000001000000000000;
                prev_state = State6_3;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State7_3)
            begin
                // Must create 5/16*Vdd
                Q = 30'b111000011000000000010000000000;
                prev_state = State6_5;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State7_3)
            begin
                // Must create 7/16*Vdd
                Q = 30'b110000011000000000011000000000;
                prev_state = State6_7;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State7_5)
            begin
                // Must create 9/16*Vdd
                Q = 30'b110011000000000000000011000000;
                prev_state = State6_9;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State7_5)
            begin
                // Must create 11/16*Vdd
                Q = 30'b110010000000000001000011000000;
                prev_state = State6_11;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State7_7)
            begin
                // Must create 13/16*Vdd
                Q = 30'b101000000000000000001111000000;
                prev_state = State6_13;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State7_7)
            begin
                // Must create 15/16*Vdd
                Q = 30'b010000000000000000001110000000;
                prev_state = State6_15;
            end
    end
  State5:
    begin
        next_state = State4;
        data_clk = 1'b1;
        get_comp = 1'b1;
        if (comp_reg == 1'b0 && prev_state_reg == State6_1)
            begin
                // Must create 1/32*Vdd
                Q = 30'b010001001100000000000000000000;
                prev_state = State5_1;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State6_1)
            begin
                // Must create 3/32*Vdd
                Q = 30'b010000001111000100000000000000;
                prev_state = State5_3;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State6_3)
            begin
                // Must create 5/32*Vdd
                Q = 30'b110001000100000000000000000000;
                prev_state = State5_5;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State6_3)
            begin
                // Must create 7/32*Vdd
                Q = 30'b100010000111000000100000000000;
                prev_state = State5_7;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State6_5)
            begin
                // Must create 9/32*Vdd
                Q = 30'b111011000100000000000000000000;
                prev_state = State5_9;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State6_5)
            begin
                // Must create 11/32*Vdd
                Q = 30'b100011000110000000001000000000;
                prev_state = State5_11;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State6_7)
            begin
                // Must create 13/32*Vdd
                Q = 30'b100000000111000000000110000000;
                prev_state = State5_13;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State6_7)
            begin
                // Must create 15/32*Vdd
                Q = 30'b100010000110000000000110000000;
                prev_state = State5_15;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State6_9)
            begin
                // Must create 17/32*Vdd
                Q = 30'b101000110000000000000000110000;
                prev_state = State5_17;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State6_9)
            begin
                // Must create 19/32*Vdd
                Q = 30'b100000110000000000000000111000;
                prev_state = State5_19;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State6_11)
            begin
                // Must create 21/32*Vdd
                Q = 30'b101101000000000000000000110000;
                prev_state = State5_21;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State6_11)
            begin
                // Must create 23/32*Vdd
                Q = 30'b111110000000000000000000100000;
                prev_state = State5_23;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State6_13)
            begin
                // Must create 25/32*Vdd
                Q = 30'b100100000000000000010000111000;
                prev_state = State5_25;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State6_13)
            begin
                // Must create 27/32*Vdd
                Q = 30'b111000000000000000000000100000;
                prev_state = State5_27;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State6_15)
            begin
                // Must create 29/32*Vdd
                Q = 30'b010000000000000100000001111000;
                prev_state = State5_29;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State6_15)
            begin
                // Must create 31/32*Vdd
                Q = 30'b010000000000000000001001100000;
                prev_state = State5_31;
            end
    end
  State4:
    begin
        next_state = State3;
        data_clk = 1'b1;
        get_comp = 1'b1;
        if (comp_reg == 1'b0 && prev_state_reg == State5_1)
            begin
                // Must create 1/64*Vdd
                Q = 30'b010000000010000000000000000000;
                prev_state = State4_1;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_1)
            begin
                // Must create 3/64*Vdd
                Q = 30'b011000000011110000000000000000;
                prev_state = State4_3;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_3)
            begin
                // Must create 5/64*Vdd
                Q = 30'b010000001111100000000000000000;
                prev_state = State4_5;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_3)
            begin
                // Must create 7/64*Vdd
                Q = 30'b011001101100000000000000000000;
                prev_state = State4_7;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_5)
            begin
                // Must create 9/64*Vdd
                Q = 30'b110001110010000000000000000000;
                prev_state = State4_9;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_5)
            begin
                // Must create 11/64*Vdd
                Q = 30'b100000110011000100000000000000;
                prev_state = State4_11;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_7)
            begin
                // Must create 13/64*Vdd
                Q = 30'b111000000000110100000000000000;
                prev_state = State4_13;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_7)
            begin
                // Must create 15/64*Vdd
                Q = 30'b100010000000100100000000000000;
                prev_state = State4_15;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_9)
            begin
                // Must create 17/64*Vdd
                Q = 30'b100000111010000000010000000000;
                prev_state = State4_17;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_9)
            begin
                // Must create 19/64*Vdd
                Q = 30'b111100110000000000000000000000;
                prev_state = State4_19;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_11)
            begin
                // Must create 21/64*Vdd
                Q = 30'b111000000001100000000100000000;
                prev_state = State4_21;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_11)
            begin
                // Must create 23/64*Vdd
                Q = 30'b110000000001100100000100000000;
                prev_state = State4_23;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_13)
            begin
                // Must create 25/64*Vdd
                Q = 30'b100011100110000000000000000000;
                prev_state = State4_25;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_13)
            begin
                // Must create 27/64*Vdd
                Q = 30'b110000011110000000000000000000;
                prev_state = State4_27;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_15)
            begin
                // Must create 29/64*Vdd
                Q = 30'b110010011100000000000000000000;
                prev_state = State4_29;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_15)
            begin
                // Must create 31/64*Vdd
                Q = 30'b110000000001100000000001100000;
                prev_state = State4_31;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_17)
            begin
                // Must create 33/64*Vdd
                Q = 30'b110000001100000000000000001100;
                prev_state = State4_33;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_17)
            begin
                // Must create 35/64*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State4_35;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_19)
            begin
                // Must create 37/64*Vdd
                Q = 30'b110011110000000000000000000000;
                prev_state = State4_37;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_19)
            begin
                // Must create 39/64*Vdd
                Q = 30'b101100110000000000010000000000;
                prev_state = State4_39;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_21)
            begin
                // Must create 41/64*Vdd
                Q = 30'b110000100000000100000000001100;
                prev_state = State4_41;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_21)
            begin
                // Must create 43/64*Vdd
                Q = 30'b110010100000000000000000001100;
                prev_state = State4_43;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_23)
            begin
                // Must create 45/64*Vdd
                Q = 30'b111000000000000001110000000000;
                prev_state = State4_45;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_23)
            begin
                // Must create 47/64*Vdd
                Q = 30'b100000000000000001010011010000;
                prev_state = State4_47;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_25)
            begin
                // Must create 49/64*Vdd
                Q = 30'b100100000000000100000000000100;
                prev_state = State4_49;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_25)
            begin
                // Must create 51/64*Vdd
                Q = 30'b110000000000000101000000000110;
                prev_state = State4_51;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_27)
            begin
                // Must create 53/64*Vdd
                Q = 30'b100000000000000100001100011000;
                prev_state = State4_53;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_27)
            begin
                // Must create 55/64*Vdd
                Q = 30'b111000000000000000001100010000;
                prev_state = State4_55;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_29)
            begin
                // Must create 57/64*Vdd
                Q = 30'b010000000000000101001101000000;
                prev_state = State4_57;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_29)
            begin
                // Must create 59/64*Vdd
                Q = 30'b010000000000000100000001110100;
                prev_state = State4_59;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State5_31)
            begin
                // Must create 61/64*Vdd
                Q = 30'b010000000000000001000000011110;
                prev_state = State4_61;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State5_31)
            begin
                // Must create 63/64*Vdd
                Q = 30'b010000000000000000000000010000;
                prev_state = State4_63;
            end
    end
  State3:
    begin
        next_state = State2;
        data_clk = 1'b1;
        get_comp = 1'b1;
        if (comp_reg == 1'b0 && prev_state_reg == State4_1)
            begin
                // Must create 1/128*Vdd
                Q = 30'b010000000001000000000000000000;
                prev_state = State3_1;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_1)
            begin
                // Must create 3/128*Vdd
                Q = 30'b010000100011000000000000000000;
                prev_state = State3_3;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_3)
            begin
                // Must create 5/128*Vdd
                Q = 30'b011000000011101000000000000000;
                prev_state = State3_5;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_3)
            begin
                // Must create 7/128*Vdd
                Q = 30'b111001001010000000000000000000;
                prev_state = State3_7;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_5)
            begin
                // Must create 9/128*Vdd
                Q = 30'b110001001100010000000000000000;
                prev_state = State3_9;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_5)
            begin
                // Must create 11/128*Vdd
                Q = 30'b110000001111000000000000000000;
                prev_state = State3_11;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_7)
            begin
                // Must create 13/128*Vdd
                Q = 30'b011001111000000000000000000000;
                prev_state = State3_13;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_7)
            begin
                // Must create 15/128*Vdd
                Q = 30'b010100010011000100000000000000;
                prev_state = State3_15;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_9)
            begin
                // Must create 17/128*Vdd
                Q = 30'b110001001001000001000000000000;
                prev_state = State3_17;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_9)
            begin
                // Must create 19/128*Vdd
                Q = 30'b101000000001110100000000000000;
                prev_state = State3_19;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_11)
            begin
                // Must create 21/128*Vdd
                Q = 30'b100010110011000000000000000000;
                prev_state = State3_21;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_11)
            begin
                // Must create 23/128*Vdd
                Q = 30'b111001110000000000000000000000;
                prev_state = State3_23;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_13)
            begin
                // Must create 25/128*Vdd
                Q = 30'b110001100000000000000000000000;
                prev_state = State3_25;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_13)
            begin
                // Must create 27/128*Vdd
                Q = 30'b111010000110000000000000000000;
                prev_state = State3_27;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_15)
            begin
                // Must create 29/128*Vdd
                Q = 30'b100010000111100000000000000000;
                prev_state = State3_29;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_15)
            begin
                // Must create 31/128*Vdd
                Q = 30'b100010000000010010000000000000;
                prev_state = State3_31;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_17)
            begin
                // Must create 33/128*Vdd
                Q = 30'b100000110001000001100000000000;
                prev_state = State3_33;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_17)
            begin
                // Must create 35/128*Vdd
                Q = 30'b111010110000000000000000000000;
                prev_state = State3_35;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_19)
            begin
                // Must create 37/128*Vdd
                Q = 30'b000010000010000101000000000000;
                prev_state = State3_37;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_19)
            begin
                // Must create 39/128*Vdd
                Q = 30'b111011000000000001000000000000;
                prev_state = State3_39;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_21)
            begin
                // Must create 41/128*Vdd
                Q = 30'b100110000000011000000010000000;
                prev_state = State3_41;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_21)
            begin
                // Must create 43/128*Vdd
                Q = 30'b100011000000011000000010000000;
                prev_state = State3_43;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_23)
            begin
                // Must create 45/128*Vdd
                Q = 30'b110011000101000000000000000000;
                prev_state = State3_45;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_23)
            begin
                // Must create 47/128*Vdd
                Q = 30'b100010000000011010000010000000;
                prev_state = State3_47;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_25)
            begin
                // Must create 49/128*Vdd
                Q = 30'b111000000001000000000110000000;
                prev_state = State3_49;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_25)
            begin
                // Must create 51/128*Vdd
                Q = 30'b100000000000111000000001100000;
                prev_state = State3_51;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_27)
            begin
                // Must create 53/128*Vdd
                Q = 30'b110000010001000000000110000000;
                prev_state = State3_53;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_27)
            begin
                // Must create 55/128*Vdd
                Q = 30'b100011000001100000000001000000;
                prev_state = State3_55;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_29)
            begin
                // Must create 57/128*Vdd
                Q = 30'b110011000010000000000100000000;
                prev_state = State3_57;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_29)
            begin
                // Must create 59/128*Vdd
                Q = 30'b110010000010000000000110000000;
                prev_state = State3_59;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_31)
            begin
                // Must create 61/128*Vdd
                Q = 30'b110010000111000000000000000000;
                prev_state = State3_61;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_31)
            begin
                // Must create 63/128*Vdd
                Q = 30'b100010000000011000000000011000;
                prev_state = State3_63;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_33)
            begin
                // Must create 65/128*Vdd
                Q = 30'b101000000011000000000000000011;
                prev_state = State3_65;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_33)
            begin
                // Must create 67/128*Vdd
                Q = 30'b111000111000000000000000000000;
                prev_state = State3_67;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_35)
            begin
                // Must create 69/128*Vdd
                Q = 30'b111000010000000000000000110000;
                prev_state = State3_69;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_35)
            begin
                // Must create 71/128*Vdd
                Q = 30'b111100010000000000000000100000;
                prev_state = State3_71;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_37)
            begin
                // Must create 73/128*Vdd
                Q = 30'b101100001000000000000000100100;
                prev_state = State3_73;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_37)
            begin
                // Must create 75/128*Vdd
                Q = 30'b110010000000000000000000111000;
                prev_state = State3_75;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_39)
            begin
                // Must create 77/128*Vdd
                Q = 30'b100000001100000000000000000111;
                prev_state = State3_77;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_39)
            begin
                // Must create 79/128*Vdd
                Q = 30'b110000000000000001000000111000;
                prev_state = State3_79;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_41)
            begin
                // Must create 81/128*Vdd
                Q = 30'b101000010000000010000000000011;
                prev_state = State3_81;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_41)
            begin
                // Must create 83/128*Vdd
                Q = 30'b111101100000000000000000000000;
                prev_state = State3_83;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_43)
            begin
                // Must create 85/128*Vdd
                Q = 30'b101100010000000000000000000011;
                prev_state = State3_85;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_43)
            begin
                // Must create 87/128*Vdd
                Q = 30'b101000010000000000100000000011;
                prev_state = State3_87;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_45)
            begin
                // Must create 89/128*Vdd
                Q = 30'b111110000000000000001000000000;
                prev_state = State3_89;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_45)
            begin
                // Must create 91/128*Vdd
                Q = 30'b000100000000000100001000010000;
                prev_state = State3_91;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_47)
            begin
                // Must create 93/128*Vdd
                Q = 30'b111100000000000001010000000000;
                prev_state = State3_93;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_47)
            begin
                // Must create 95/128*Vdd
                Q = 30'b100000000000000001011100001000;
                prev_state = State3_95;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_49)
            begin
                // Must create 97/128*Vdd
                Q = 30'b100100000000000010000000000010;
                prev_state = State3_97;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_49)
            begin
                // Must create 99/128*Vdd
                Q = 30'b100100000000000100010000110000;
                prev_state = State3_99;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_51)
            begin
                // Must create 101/128*Vdd
                Q = 30'b110100000000000100010000100000;
                prev_state = State3_101;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_51)
            begin
                // Must create 103/128*Vdd
                Q = 30'b111000000000000000001000000000;
                prev_state = State3_103;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_53)
            begin
                // Must create 105/128*Vdd
                Q = 30'b111000000000000101001000000000;
                prev_state = State3_105;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_53)
            begin
                // Must create 107/128*Vdd
                Q = 30'b100000000000000100011100010000;
                prev_state = State3_107;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_55)
            begin
                // Must create 109/128*Vdd
                Q = 30'b100000000000000101000000001110;
                prev_state = State3_109;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_55)
            begin
                // Must create 111/128*Vdd
                Q = 30'b111000000000000000000011001000;
                prev_state = State3_111;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_57)
            begin
                // Must create 113/128*Vdd
                Q = 30'b010000000000000000100010111000;
                prev_state = State3_113;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_57)
            begin
                // Must create 115/128*Vdd
                Q = 30'b010000000000000101001110000000;
                prev_state = State3_115;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_59)
            begin
                // Must create 117/128*Vdd
                Q = 30'b110000000000000100000001110000;
                prev_state = State3_117;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_59)
            begin
                // Must create 119/128*Vdd
                Q = 30'b110000000000000100001001000010;
                prev_state = State3_119;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_61)
            begin
                // Must create 121/128*Vdd
                Q = 30'b110000000000000001001001010000;
                prev_state = State3_121;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_61)
            begin
                // Must create 123/128*Vdd
                Q = 30'b010000000000000001000000011101;
                prev_state = State3_123;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State4_63)
            begin
                // Must create 125/128*Vdd
                Q = 30'b010000000000000000000100011000;
                prev_state = State3_125;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State4_63)
            begin
                // Must create 127/128*Vdd
                Q = 30'b010000000000000000000000001000;
                prev_state = State3_127;
            end
    end
  State2:
    begin
        next_state = State1;
        data_clk = 1'b1;
        get_comp = 1'b1;
        if (comp_reg == 1'b0 && prev_state_reg == State3_1)
            begin
                // Must create 1/256*Vdd
                Q = 30'b010000000000100000000000000000;
                prev_state = State2_1;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_1)
            begin
                // Must create 3/256*Vdd
                Q = 30'b010001000001100000000000000000;
                prev_state = State2_3;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_3)
            begin
                // Must create 5/256*Vdd
                Q = 30'b010001100000100000000000000000;
                prev_state = State2_5;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_3)
            begin
                // Must create 7/256*Vdd
                Q = 30'b010001101000000000000000000000;
                prev_state = State2_7;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_5)
            begin
                // Must create 9/256*Vdd
                Q = 30'b010001000000000000000000000000;
                prev_state = State2_9;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_5)
            begin
                // Must create 11/256*Vdd
                Q = 30'b011000100011100000000000000000;
                prev_state = State2_11;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_7)
            begin
                // Must create 13/256*Vdd
                Q = 30'b111001001100000000000000000000;
                prev_state = State2_13;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_7)
            begin
                // Must create 15/256*Vdd
                Q = 30'b100010000101110000000000000000;
                prev_state = State2_15;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_9)
            begin
                // Must create 17/256*Vdd
                Q = 30'b100000000011101100000000000000;
                prev_state = State2_17;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_9)
            begin
                // Must create 19/256*Vdd
                Q = 30'b110001001100000100000000000000;
                prev_state = State2_19;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_11)
            begin
                // Must create 21/256*Vdd
                Q = 30'b110001001110000000000000000000;
                prev_state = State2_21;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_11)
            begin
                // Must create 23/256*Vdd
                Q = 30'b101001100000110000000000000000;
                prev_state = State2_23;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_13)
            begin
                // Must create 25/256*Vdd
                Q = 30'b110100000100110000000000000000;
                prev_state = State2_25;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_13)
            begin
                // Must create 27/256*Vdd
                Q = 30'b111001110000000000000000000000;
                prev_state = State2_27;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_15)
            begin
                // Must create 29/256*Vdd
                Q = 30'b011101110000000000000000000000;
                prev_state = State2_29;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_15)
            begin
                // Must create 31/256*Vdd
                Q = 30'b011000000000111010000000000000;
                prev_state = State2_31;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_17)
            begin
                // Must create 33/256*Vdd
                Q = 30'b111000000000100000000000000000;
                prev_state = State2_33;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_17)
            begin
                // Must create 35/256*Vdd
                Q = 30'b110001001101000000000000000000;
                prev_state = State2_35;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_19)
            begin
                // Must create 37/256*Vdd
                Q = 30'b111001100001000000000000000000;
                prev_state = State2_37;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_19)
            begin
                // Must create 39/256*Vdd
                Q = 30'b111001001001000000000000000000;
                prev_state = State2_39;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_21)
            begin
                // Must create 41/256*Vdd
                Q = 30'b101000001000100101000000000000;
                prev_state = State2_41;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_21)
            begin
                // Must create 43/256*Vdd
                Q = 30'b100010111010000000000000000000;
                prev_state = State2_43;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_23)
            begin
                // Must create 45/256*Vdd
                Q = 30'b111000000011000100000000000000;
                prev_state = State2_45;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_23)
            begin
                // Must create 47/256*Vdd
                Q = 30'b100100000111000100000000000000;
                prev_state = State2_47;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_25)
            begin
                // Must create 49/256*Vdd
                Q = 30'b100000010000000000000000000000;
                prev_state = State2_49;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_25)
            begin
                // Must create 51/256*Vdd
                Q = 30'b111001000000110000000000000000;
                prev_state = State2_51;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_27)
            begin
                // Must create 53/256*Vdd
                Q = 30'b111000000000110100000000000000;
                prev_state = State2_53;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_27)
            begin
                // Must create 55/256*Vdd
                Q = 30'b111100000000110000000000000000;
                prev_state = State2_55;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_29)
            begin
                // Must create 57/256*Vdd
                Q = 30'b110011000100000000100000000000;
                prev_state = State2_57;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_29)
            begin
                // Must create 59/256*Vdd
                Q = 30'b110010000111000000000000000000;
                prev_state = State2_59;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_31)
            begin
                // Must create 61/256*Vdd
                Q = 30'b110010000100110000000000000000;
                prev_state = State2_61;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_31)
            begin
                // Must create 63/256*Vdd
                Q = 30'b110000000000000000000000000000;
                prev_state = State2_63;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_33)
            begin
                // Must create 65/256*Vdd
                Q = 30'b100000100000100100000000000000;
                prev_state = State2_65;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_33)
            begin
                // Must create 67/256*Vdd
                Q = 30'b100000111010000000010000000000;
                prev_state = State2_67;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_35)
            begin
                // Must create 69/256*Vdd
                Q = 30'b111000001010000000010000000000;
                prev_state = State2_69;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_35)
            begin
                // Must create 71/256*Vdd
                Q = 30'b100100001001000101000000000000;
                prev_state = State2_71;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_37)
            begin
                // Must create 73/256*Vdd
                Q = 30'b100010001001000010010000000000;
                prev_state = State2_73;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_37)
            begin
                // Must create 75/256*Vdd
                Q = 30'b111010000010000100000000000000;
                prev_state = State2_75;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_39)
            begin
                // Must create 77/256*Vdd
                Q = 30'b111100110000000000000000000000;
                prev_state = State2_77;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_39)
            begin
                // Must create 79/256*Vdd
                Q = 30'b100100110100000000100000000000;
                prev_state = State2_79;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_41)
            begin
                // Must create 81/256*Vdd
                Q = 30'b100000010000000000000000000000;
                prev_state = State2_81;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_41)
            begin
                // Must create 83/256*Vdd
                Q = 30'b111110000001000000000000000000;
                prev_state = State2_83;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_43)
            begin
                // Must create 85/256*Vdd
                Q = 30'b111011000001000000000000000000;
                prev_state = State2_85;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_43)
            begin
                // Must create 87/256*Vdd
                Q = 30'b100011000110000000001000000000;
                prev_state = State2_87;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_45)
            begin
                // Must create 89/256*Vdd
                Q = 30'b111010000000100100000000000000;
                prev_state = State2_89;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_45)
            begin
                // Must create 91/256*Vdd
                Q = 30'b110010000000100100000100000000;
                prev_state = State2_91;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_47)
            begin
                // Must create 93/256*Vdd
                Q = 30'b110010000001110000000000000000;
                prev_state = State2_93;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_47)
            begin
                // Must create 95/256*Vdd
                Q = 30'b100000100000000000000000000000;
                prev_state = State2_95;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_49)
            begin
                // Must create 97/256*Vdd
                Q = 30'b111100011000000000000000000000;
                prev_state = State2_97;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_49)
            begin
                // Must create 99/256*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State2_99;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_51)
            begin
                // Must create 101/256*Vdd
                Q = 30'b100011100000110000000000000000;
                prev_state = State2_101;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_51)
            begin
                // Must create 103/256*Vdd
                Q = 30'b100000000001110000000110000000;
                prev_state = State2_103;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_53)
            begin
                // Must create 105/256*Vdd
                Q = 30'b110010011100000000000000000000;
                prev_state = State2_105;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_53)
            begin
                // Must create 107/256*Vdd
                Q = 30'b110000011110000000000000000000;
                prev_state = State2_107;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_55)
            begin
                // Must create 109/256*Vdd
                Q = 30'b110011011000000000000000000000;
                prev_state = State2_109;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_55)
            begin
                // Must create 111/256*Vdd
                Q = 30'b110000100000010001000000100000;
                prev_state = State2_111;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_57)
            begin
                // Must create 113/256*Vdd
                Q = 30'b100000111100000000000010000000;
                prev_state = State2_113;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_57)
            begin
                // Must create 115/256*Vdd
                Q = 30'b110010011100000000000000000000;
                prev_state = State2_115;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_59)
            begin
                // Must create 117/256*Vdd
                Q = 30'b110010011100000000000000000000;
                prev_state = State2_117;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_59)
            begin
                // Must create 119/256*Vdd
                Q = 30'b100000010001000000011001000000;
                prev_state = State2_119;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_61)
            begin
                // Must create 121/256*Vdd
                Q = 30'b110010010000100000000001000000;
                prev_state = State2_121;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_61)
            begin
                // Must create 123/256*Vdd
                Q = 30'b110010000000100000000001100000;
                prev_state = State2_123;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_63)
            begin
                // Must create 125/256*Vdd
                Q = 30'b110010000001110000000000000000;
                prev_state = State2_125;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_63)
            begin
                // Must create 127/256*Vdd
                Q = 30'b111001100000000000000000000100;
                prev_state = State2_127;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_65)
            begin
                // Must create 129/256*Vdd
                Q = 30'b110100000000100001010000000000;
                prev_state = State2_129;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_65)
            begin
                // Must create 131/256*Vdd
                Q = 30'b111000001110000000000000000000;
                prev_state = State2_131;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_67)
            begin
                // Must create 133/256*Vdd
                Q = 30'b111000000100000000000000001100;
                prev_state = State2_133;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_67)
            begin
                // Must create 135/256*Vdd
                Q = 30'b111010000100000000000000001000;
                prev_state = State2_135;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_69)
            begin
                // Must create 137/256*Vdd
                Q = 30'b100010001000000000000011001000;
                prev_state = State2_137;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_69)
            begin
                // Must create 139/256*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State2_139;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_71)
            begin
                // Must create 141/256*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State2_141;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_71)
            begin
                // Must create 143/256*Vdd
                Q = 30'b100011100000000000010000010000;
                prev_state = State2_143;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_73)
            begin
                // Must create 145/256*Vdd
                Q = 30'b110000000100000000011000000010;
                prev_state = State2_145;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_73)
            begin
                // Must create 147/256*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State2_147;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_75)
            begin
                // Must create 149/256*Vdd
                Q = 30'b110011110000000000000000000000;
                prev_state = State2_149;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_75)
            begin
                // Must create 151/256*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State2_151;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_77)
            begin
                // Must create 153/256*Vdd
                Q = 30'b100000001100000000000000111000;
                prev_state = State2_153;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_77)
            begin
                // Must create 155/256*Vdd
                Q = 30'b101100101100000000000000000000;
                prev_state = State2_155;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_79)
            begin
                // Must create 157/256*Vdd
                Q = 30'b111100100000000001000000000000;
                prev_state = State2_157;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_79)
            begin
                // Must create 159/256*Vdd
                Q = 30'b110011000000000001100000000000;
                prev_state = State2_159;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_81)
            begin
                // Must create 161/256*Vdd
                Q = 30'b100000000000000000010000000000;
                prev_state = State2_161;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_81)
            begin
                // Must create 163/256*Vdd
                Q = 30'b111000110000000100000000000000;
                prev_state = State2_163;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_83)
            begin
                // Must create 165/256*Vdd
                Q = 30'b111000000000000100000000001100;
                prev_state = State2_165;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_83)
            begin
                // Must create 167/256*Vdd
                Q = 30'b111010000000000100000000001000;
                prev_state = State2_167;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_85)
            begin
                // Must create 169/256*Vdd
                Q = 30'b101101000000000000000000110000;
                prev_state = State2_169;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_85)
            begin
                // Must create 171/256*Vdd
                Q = 30'b111110100000000000000000000000;
                prev_state = State2_171;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_87)
            begin
                // Must create 173/256*Vdd
                Q = 30'b111010110000000000000000000000;
                prev_state = State2_173;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_87)
            begin
                // Must create 175/256*Vdd
                Q = 30'b100000000000000001000000000000;
                prev_state = State2_175;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_89)
            begin
                // Must create 177/256*Vdd
                Q = 30'b100000000000000001110100100000;
                prev_state = State2_177;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_89)
            begin
                // Must create 179/256*Vdd
                Q = 30'b111000000000000001110000000000;
                prev_state = State2_179;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_91)
            begin
                // Must create 181/256*Vdd
                Q = 30'b111100000000000100001000000000;
                prev_state = State2_181;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_91)
            begin
                // Must create 183/256*Vdd
                Q = 30'b100100000000000010000011001000;
                prev_state = State2_183;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_93)
            begin
                // Must create 185/256*Vdd
                Q = 30'b100000000000000100101010001000;
                prev_state = State2_185;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_93)
            begin
                // Must create 187/256*Vdd
                Q = 30'b111000000000000000000011010000;
                prev_state = State2_187;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_95)
            begin
                // Must create 189/256*Vdd
                Q = 30'b100000000000000001010011010000;
                prev_state = State2_189;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_95)
            begin
                // Must create 191/256*Vdd
                Q = 30'b100000000000000101000000000100;
                prev_state = State2_191;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_97)
            begin
                // Must create 193/256*Vdd
                Q = 30'b110000000000000000000000000000;
                prev_state = State2_193;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_97)
            begin
                // Must create 195/256*Vdd
                Q = 30'b110100000000000110010000000000;
                prev_state = State2_195;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_99)
            begin
                // Must create 197/256*Vdd
                Q = 30'b110100000000000100010000100000;
                prev_state = State2_197;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_99)
            begin
                // Must create 199/256*Vdd
                Q = 30'b111100000000000100000000001000;
                prev_state = State2_199;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_101)
            begin
                // Must create 201/256*Vdd
                Q = 30'b110100000000000001100000000100;
                prev_state = State2_201;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_101)
            begin
                // Must create 203/256*Vdd
                Q = 30'b110100000000000001000000000110;
                prev_state = State2_203;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_103)
            begin
                // Must create 205/256*Vdd
                Q = 30'b111000000000000101000000000100;
                prev_state = State2_205;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_103)
            begin
                // Must create 207/256*Vdd
                Q = 30'b100000000000000000000100000000;
                prev_state = State2_207;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_105)
            begin
                // Must create 209/256*Vdd
                Q = 30'b100000000000000000100100111000;
                prev_state = State2_209;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_105)
            begin
                // Must create 211/256*Vdd
                Q = 30'b111000000000000000000100011000;
                prev_state = State2_211;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_107)
            begin
                // Must create 213/256*Vdd
                Q = 30'b100000000000000100011110000000;
                prev_state = State2_213;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_107)
            begin
                // Must create 215/256*Vdd
                Q = 30'b100000000000000001000011001100;
                prev_state = State2_215;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_109)
            begin
                // Must create 217/256*Vdd
                Q = 30'b111000000000000101000010000000;
                prev_state = State2_217;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_109)
            begin
                // Must create 219/256*Vdd
                Q = 30'b111000000000000101001000000000;
                prev_state = State2_219;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_111)
            begin
                // Must create 221/256*Vdd
                Q = 30'b111000000000000000000011100000;
                prev_state = State2_221;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_111)
            begin
                // Must create 223/256*Vdd
                Q = 30'b110000000000000001000000000100;
                prev_state = State2_223;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_113)
            begin
                // Must create 225/256*Vdd
                Q = 30'b010000000000000110000000000111;
                prev_state = State2_225;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_113)
            begin
                // Must create 227/256*Vdd
                Q = 30'b010000000000000101101010000000;
                prev_state = State2_227;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_115)
            begin
                // Must create 229/256*Vdd
                Q = 30'b110000000000000101001100000000;
                prev_state = State2_229;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_115)
            begin
                // Must create 231/256*Vdd
                Q = 30'b110000000000000000100001000110;
                prev_state = State2_231;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_117)
            begin
                // Must create 233/256*Vdd
                Q = 30'b100000000000000001001100000110;
                prev_state = State2_233;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_117)
            begin
                // Must create 235/256*Vdd
                Q = 30'b110000000000000100001001100000;
                prev_state = State2_235;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_119)
            begin
                // Must create 237/256*Vdd
                Q = 30'b110000000000000100001001001000;
                prev_state = State2_237;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_119)
            begin
                // Must create 239/256*Vdd
                Q = 30'b100000000000000000000000111101;
                prev_state = State2_239;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_121)
            begin
                // Must create 241/256*Vdd
                Q = 30'b100000000000000000010000101110;
                prev_state = State2_241;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_121)
            begin
                // Must create 243/256*Vdd
                Q = 30'b110000000000000001001001100000;
                prev_state = State2_243;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_123)
            begin
                // Must create 245/256*Vdd
                Q = 30'b010000000000000001000100011100;
                prev_state = State2_245;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_123)
            begin
                // Must create 247/256*Vdd
                Q = 30'b010000000000000000001000000000;
                prev_state = State2_247;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_125)
            begin
                // Must create 249/256*Vdd
                Q = 30'b010000000000000000001101000000;
                prev_state = State2_249;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_125)
            begin
                // Must create 251/256*Vdd
                Q = 30'b010000000000000000001100000100;
                prev_state = State2_251;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State3_127)
            begin
                // Must create 253/256*Vdd
                Q = 30'b010000000000000000001000001100;
                prev_state = State2_253;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State3_127)
            begin
                // Must create 255/256*Vdd
                Q = 30'b010000000000000000000000000100;
                prev_state = State2_255;
            end
    end
  State1:
    begin
        next_state = State0;
        data_clk = 1'b1;
        get_comp = 1'b1;
        if (comp_reg == 1'b0 && prev_state_reg == State2_1)
            begin
                // Must create 1/512*Vdd
                Q = 30'b010000000000010000000000000000;
                prev_state = State1_1;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_1)
            begin
                // Must create 3/512*Vdd
                Q = 30'b010000000010110000000000000000;
                prev_state = State1_3;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_3)
            begin
                // Must create 5/512*Vdd
                Q = 30'b010001000010010000000000000000;
                prev_state = State1_5;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_3)
            begin
                // Must create 7/512*Vdd
                Q = 30'b010001001011010000000000000000;
                prev_state = State1_7;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_5)
            begin
                // Must create 9/512*Vdd
                Q = 30'b010001100011010000000000000000;
                prev_state = State1_9;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_5)
            begin
                // Must create 11/512*Vdd
                Q = 30'b010000010011011000000000000000;
                prev_state = State1_11;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_7)
            begin
                // Must create 13/512*Vdd
                Q = 30'b010001000011000000000000000000;
                prev_state = State1_13;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_7)
            begin
                // Must create 15/512*Vdd
                Q = 30'b110000000010111000000000000000;
                prev_state = State1_15;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_9)
            begin
                // Must create 17/512*Vdd
                Q = 30'b010000001000000000000000000000;
                prev_state = State1_17;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_9)
            begin
                // Must create 19/512*Vdd
                Q = 30'b011000001011100000000000000000;
                prev_state = State1_19;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_11)
            begin
                // Must create 21/512*Vdd
                Q = 30'b011001100011000000000000000000;
                prev_state = State1_21;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_11)
            begin
                // Must create 23/512*Vdd
                Q = 30'b011001010000000000000000000000;
                prev_state = State1_23;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_13)
            begin
                // Must create 25/512*Vdd
                Q = 30'b110000000001100000000000000000;
                prev_state = State1_25;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_13)
            begin
                // Must create 27/512*Vdd
                Q = 30'b111001101000000000000000000000;
                prev_state = State1_27;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_15)
            begin
                // Must create 29/512*Vdd
                Q = 30'b111011000100000000000000000000;
                prev_state = State1_29;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_15)
            begin
                // Must create 31/512*Vdd
                Q = 30'b100000100000000000000000000000;
                prev_state = State1_31;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_17)
            begin
                // Must create 33/512*Vdd
                Q = 30'b100000100000000000000000000000;
                prev_state = State1_33;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_17)
            begin
                // Must create 35/512*Vdd
                Q = 30'b110001001011000000000000000000;
                prev_state = State1_35;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_19)
            begin
                // Must create 37/512*Vdd
                Q = 30'b110001101100000000000000000000;
                prev_state = State1_37;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_19)
            begin
                // Must create 39/512*Vdd
                Q = 30'b110000000011000000000000000000;
                prev_state = State1_39;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_21)
            begin
                // Must create 41/512*Vdd
                Q = 30'b110001100000100100000000000000;
                prev_state = State1_41;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_21)
            begin
                // Must create 43/512*Vdd
                Q = 30'b110001001100000100000000000000;
                prev_state = State1_43;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_23)
            begin
                // Must create 45/512*Vdd
                Q = 30'b111001001100000000000000000000;
                prev_state = State1_45;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_23)
            begin
                // Must create 47/512*Vdd
                Q = 30'b101010010000000000000000000000;
                prev_state = State1_47;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_25)
            begin
                // Must create 49/512*Vdd
                Q = 30'b110000000011000000000000000000;
                prev_state = State1_49;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_25)
            begin
                // Must create 51/512*Vdd
                Q = 30'b111101100000000000000000000000;
                prev_state = State1_51;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_27)
            begin
                // Must create 53/512*Vdd
                Q = 30'b111001100010000000000000000000;
                prev_state = State1_53;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_27)
            begin
                // Must create 55/512*Vdd
                Q = 30'b111010000110000000000000000000;
                prev_state = State1_55;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_29)
            begin
                // Must create 57/512*Vdd
                Q = 30'b010000001000000000000000000000;
                prev_state = State1_57;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_29)
            begin
                // Must create 59/512*Vdd
                Q = 30'b011100000011000100000000000000;
                prev_state = State1_59;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_31)
            begin
                // Must create 61/512*Vdd
                Q = 30'b011100010010100000000000000000;
                prev_state = State1_61;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_31)
            begin
                // Must create 63/512*Vdd
                Q = 30'b110000000000000000000000000000;
                prev_state = State1_63;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_33)
            begin
                // Must create 65/512*Vdd
                Q = 30'b110100000000010000000000000000;
                prev_state = State1_65;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_33)
            begin
                // Must create 67/512*Vdd
                Q = 30'b111001001001000000000000000000;
                prev_state = State1_67;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_35)
            begin
                // Must create 69/512*Vdd
                Q = 30'b110011001100000000000000000000;
                prev_state = State1_69;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_35)
            begin
                // Must create 71/512*Vdd
                Q = 30'b110000110000000000000000000000;
                prev_state = State1_71;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_37)
            begin
                // Must create 73/512*Vdd
                Q = 30'b111010000000110000000000000000;
                prev_state = State1_73;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_37)
            begin
                // Must create 75/512*Vdd
                Q = 30'b111000000000110100000000000000;
                prev_state = State1_75;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_39)
            begin
                // Must create 77/512*Vdd
                Q = 30'b111000000000110100000000000000;
                prev_state = State1_77;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_39)
            begin
                // Must create 79/512*Vdd
                Q = 30'b100000100000110101000000000000;
                prev_state = State1_79;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_41)
            begin
                // Must create 81/512*Vdd
                Q = 30'b111001000000000000000000000000;
                prev_state = State1_81;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_41)
            begin
                // Must create 83/512*Vdd
                Q = 30'b101010111000000000000000000000;
                prev_state = State1_83;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_43)
            begin
                // Must create 85/512*Vdd
                Q = 30'b110010111000000000000000000000;
                prev_state = State1_85;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_43)
            begin
                // Must create 87/512*Vdd
                Q = 30'b101100000001100001000000000000;
                prev_state = State1_87;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_45)
            begin
                // Must create 89/512*Vdd
                Q = 30'b111001100100000000000000000000;
                prev_state = State1_89;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_45)
            begin
                // Must create 91/512*Vdd
                Q = 30'b111001110000000000000000000000;
                prev_state = State1_91;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_47)
            begin
                // Must create 93/512*Vdd
                Q = 30'b111101000100000000000000000000;
                prev_state = State1_93;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_47)
            begin
                // Must create 95/512*Vdd
                Q = 30'b100000001000000000000000000000;
                prev_state = State1_95;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_49)
            begin
                // Must create 97/512*Vdd
                Q = 30'b100000001000000000000000000000;
                prev_state = State1_97;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_49)
            begin
                // Must create 99/512*Vdd
                Q = 30'b111001001000000001000000000000;
                prev_state = State1_99;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_51)
            begin
                // Must create 101/512*Vdd
                Q = 30'b111001010000100000000000000000;
                prev_state = State1_101;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_51)
            begin
                // Must create 103/512*Vdd
                Q = 30'b111010010000000100000000000000;
                prev_state = State1_103;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_53)
            begin
                // Must create 105/512*Vdd
                Q = 30'b111011000100000000000000000000;
                prev_state = State1_105;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_53)
            begin
                // Must create 107/512*Vdd
                Q = 30'b111010000110000000000000000000;
                prev_state = State1_107;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_55)
            begin
                // Must create 109/512*Vdd
                Q = 30'b111010000110000000000000000000;
                prev_state = State1_109;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_55)
            begin
                // Must create 111/512*Vdd
                Q = 30'b100011100000001010000000000000;
                prev_state = State1_111;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_57)
            begin
                // Must create 113/512*Vdd
                Q = 30'b100000100011100100000000000000;
                prev_state = State1_113;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_57)
            begin
                // Must create 115/512*Vdd
                Q = 30'b110010000011100000000000000000;
                prev_state = State1_115;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_59)
            begin
                // Must create 117/512*Vdd
                Q = 30'b110010000110000000100000000000;
                prev_state = State1_117;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_59)
            begin
                // Must create 119/512*Vdd
                Q = 30'b111010000000000100100000000000;
                prev_state = State1_119;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_61)
            begin
                // Must create 121/512*Vdd
                Q = 30'b111010000010000100000000000000;
                prev_state = State1_121;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_61)
            begin
                // Must create 123/512*Vdd
                Q = 30'b111010000100100000000000000000;
                prev_state = State1_123;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_63)
            begin
                // Must create 125/512*Vdd
                Q = 30'b101110000000110000000000000000;
                prev_state = State1_125;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_63)
            begin
                // Must create 127/512*Vdd
                Q = 30'b101000000000000000000000000000;
                prev_state = State1_127;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_65)
            begin
                // Must create 129/512*Vdd
                Q = 30'b100000100000010010000000000000;
                prev_state = State1_129;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_65)
            begin
                // Must create 131/512*Vdd
                Q = 30'b100000110001100001000000000000;
                prev_state = State1_131;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_67)
            begin
                // Must create 133/512*Vdd
                Q = 30'b100000110001000001100000000000;
                prev_state = State1_133;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_67)
            begin
                // Must create 135/512*Vdd
                Q = 30'b110000110001000001000000000000;
                prev_state = State1_135;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_69)
            begin
                // Must create 137/512*Vdd
                Q = 30'b111110100000000000000000000000;
                prev_state = State1_137;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_69)
            begin
                // Must create 139/512*Vdd
                Q = 30'b111010110000000000000000000000;
                prev_state = State1_139;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_71)
            begin
                // Must create 141/512*Vdd
                Q = 30'b111110001000000000000000000000;
                prev_state = State1_141;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_71)
            begin
                // Must create 143/512*Vdd
                Q = 30'b100001000000000000000000000000;
                prev_state = State1_143;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_73)
            begin
                // Must create 145/512*Vdd
                Q = 30'b100001000000000000000000000000;
                prev_state = State1_145;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_73)
            begin
                // Must create 147/512*Vdd
                Q = 30'b100010001010000101000000000000;
                prev_state = State1_147;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_75)
            begin
                // Must create 149/512*Vdd
                Q = 30'b111011000010000000000000000000;
                prev_state = State1_149;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_75)
            begin
                // Must create 151/512*Vdd
                Q = 30'b111100110000000000000000000000;
                prev_state = State1_151;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_77)
            begin
                // Must create 153/512*Vdd
                Q = 30'b111011000100000000000000000000;
                prev_state = State1_153;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_77)
            begin
                // Must create 155/512*Vdd
                Q = 30'b111011000000000001000000000000;
                prev_state = State1_155;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_79)
            begin
                // Must create 157/512*Vdd
                Q = 30'b111110100000000000000000000000;
                prev_state = State1_157;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_79)
            begin
                // Must create 159/512*Vdd
                Q = 30'b100000001000000000000000000000;
                prev_state = State1_159;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_81)
            begin
                // Must create 161/512*Vdd
                Q = 30'b100000001000000000000000000000;
                prev_state = State1_161;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_81)
            begin
                // Must create 163/512*Vdd
                Q = 30'b100110001000011000000000000000;
                prev_state = State1_163;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_83)
            begin
                // Must create 165/512*Vdd
                Q = 30'b111000000000011000000010000000;
                prev_state = State1_165;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_83)
            begin
                // Must create 167/512*Vdd
                Q = 30'b111001000000011000000000000000;
                prev_state = State1_167;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_85)
            begin
                // Must create 169/512*Vdd
                Q = 30'b111000010000011000000000000000;
                prev_state = State1_169;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_85)
            begin
                // Must create 171/512*Vdd
                Q = 30'b111000000000011000000010000000;
                prev_state = State1_171;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_87)
            begin
                // Must create 173/512*Vdd
                Q = 30'b100011000000011000000010000000;
                prev_state = State1_173;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_87)
            begin
                // Must create 175/512*Vdd
                Q = 30'b110000100000011000000010000000;
                prev_state = State1_175;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_89)
            begin
                // Must create 177/512*Vdd
                Q = 30'b100001010101000000000100000000;
                prev_state = State1_177;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_89)
            begin
                // Must create 179/512*Vdd
                Q = 30'b111001000101000000000000000000;
                prev_state = State1_179;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_91)
            begin
                // Must create 181/512*Vdd
                Q = 30'b110011000101000000000000000000;
                prev_state = State1_181;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_91)
            begin
                // Must create 183/512*Vdd
                Q = 30'b110011100100000000000000000000;
                prev_state = State1_183;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_93)
            begin
                // Must create 185/512*Vdd
                Q = 30'b110011000000001010000000000000;
                prev_state = State1_185;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_93)
            begin
                // Must create 187/512*Vdd
                Q = 30'b110010000000001010000010000000;
                prev_state = State1_187;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_95)
            begin
                // Must create 189/512*Vdd
                Q = 30'b100010000000011011000000000000;
                prev_state = State1_189;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_95)
            begin
                // Must create 191/512*Vdd
                Q = 30'b100000000000000001000000000000;
                prev_state = State1_191;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_97)
            begin
                // Must create 193/512*Vdd
                Q = 30'b100000000001110100000001000000;
                prev_state = State1_193;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_97)
            begin
                // Must create 195/512*Vdd
                Q = 30'b111000000001000000000110000000;
                prev_state = State1_195;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_99)
            begin
                // Must create 197/512*Vdd
                Q = 30'b111000000001000000000110000000;
                prev_state = State1_197;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_99)
            begin
                // Must create 199/512*Vdd
                Q = 30'b100100011001000000010000000000;
                prev_state = State1_199;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_101)
            begin
                // Must create 201/512*Vdd
                Q = 30'b100011000000001001000001000000;
                prev_state = State1_201;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_101)
            begin
                // Must create 203/512*Vdd
                Q = 30'b100011000000001000000001100000;
                prev_state = State1_203;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_103)
            begin
                // Must create 205/512*Vdd
                Q = 30'b100000000001101000000001100000;
                prev_state = State1_205;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_103)
            begin
                // Must create 207/512*Vdd
                Q = 30'b110010000000001000000001100000;
                prev_state = State1_207;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_105)
            begin
                // Must create 209/512*Vdd
                Q = 30'b100001000011000000000110000000;
                prev_state = State1_209;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_105)
            begin
                // Must create 211/512*Vdd
                Q = 30'b110010000001000000000110000000;
                prev_state = State1_211;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_107)
            begin
                // Must create 213/512*Vdd
                Q = 30'b100010000001000000011100000000;
                prev_state = State1_213;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_107)
            begin
                // Must create 215/512*Vdd
                Q = 30'b110000010001000000010100000000;
                prev_state = State1_215;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_109)
            begin
                // Must create 217/512*Vdd
                Q = 30'b110010000001100000000100000000;
                prev_state = State1_217;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_109)
            begin
                // Must create 219/512*Vdd
                Q = 30'b110010000001100000000001000000;
                prev_state = State1_219;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_111)
            begin
                // Must create 221/512*Vdd
                Q = 30'b110011100001000000000000000000;
                prev_state = State1_221;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_111)
            begin
                // Must create 223/512*Vdd
                Q = 30'b100010011000000100000100000000;
                prev_state = State1_223;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_113)
            begin
                // Must create 225/512*Vdd
                Q = 30'b110000000001000001100001000000;
                prev_state = State1_225;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_113)
            begin
                // Must create 227/512*Vdd
                Q = 30'b110011110000000000000000000000;
                prev_state = State1_227;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_115)
            begin
                // Must create 229/512*Vdd
                Q = 30'b110011000010000000000100000000;
                prev_state = State1_229;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_115)
            begin
                // Must create 231/512*Vdd
                Q = 30'b110011000010000000000010000000;
                prev_state = State1_231;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_117)
            begin
                // Must create 233/512*Vdd
                Q = 30'b110010000010000000010100000000;
                prev_state = State1_233;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_117)
            begin
                // Must create 235/512*Vdd
                Q = 30'b100001000011000000000101000000;
                prev_state = State1_235;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_119)
            begin
                // Must create 237/512*Vdd
                Q = 30'b110010010011000000000000000000;
                prev_state = State1_237;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_119)
            begin
                // Must create 239/512*Vdd
                Q = 30'b111101000000000000000000100000;
                prev_state = State1_239;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_121)
            begin
                // Must create 241/512*Vdd
                Q = 30'b100000001111000000000000100000;
                prev_state = State1_241;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_121)
            begin
                // Must create 243/512*Vdd
                Q = 30'b110010000111000000000000000000;
                prev_state = State1_243;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_123)
            begin
                // Must create 245/512*Vdd
                Q = 30'b110010000111000000000000000000;
                prev_state = State1_245;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_123)
            begin
                // Must create 247/512*Vdd
                Q = 30'b100000000100010000000110010000;
                prev_state = State1_247;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_125)
            begin
                // Must create 249/512*Vdd
                Q = 30'b110010000100001000000000010000;
                prev_state = State1_249;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_125)
            begin
                // Must create 251/512*Vdd
                Q = 30'b110010000000001000000000011000;
                prev_state = State1_251;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_127)
            begin
                // Must create 253/512*Vdd
                Q = 30'b111010000000011000000000000000;
                prev_state = State1_253;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_127)
            begin
                // Must create 255/512*Vdd
                Q = 30'b100110000000000001100000000010;
                prev_state = State1_255;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_129)
            begin
                // Must create 257/512*Vdd
                Q = 30'b101000000000010000101100000000;
                prev_state = State1_257;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_129)
            begin
                // Must create 259/512*Vdd
                Q = 30'b111100000011000000000000000000;
                prev_state = State1_259;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_131)
            begin
                // Must create 261/512*Vdd
                Q = 30'b111000000001000000000000000011;
                prev_state = State1_261;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_131)
            begin
                // Must create 263/512*Vdd
                Q = 30'b111000100001000000000000000010;
                prev_state = State1_263;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_133)
            begin
                // Must create 265/512*Vdd
                Q = 30'b100000100010000000000000110010;
                prev_state = State1_265;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_133)
            begin
                // Must create 267/512*Vdd
                Q = 30'b111000111000000000000000000000;
                prev_state = State1_267;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_135)
            begin
                // Must create 269/512*Vdd
                Q = 30'b111000111000000000000000000000;
                prev_state = State1_269;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_135)
            begin
                // Must create 271/512*Vdd
                Q = 30'b100001111000000000000000000100;
                prev_state = State1_271;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_137)
            begin
                // Must create 273/512*Vdd
                Q = 30'b110100000100000001100000000000;
                prev_state = State1_273;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_137)
            begin
                // Must create 275/512*Vdd
                Q = 30'b111010011000000000000000000000;
                prev_state = State1_275;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_139)
            begin
                // Must create 277/512*Vdd
                Q = 30'b100100011000000000000000101000;
                prev_state = State1_277;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_139)
            begin
                // Must create 279/512*Vdd
                Q = 30'b111000010000000000000010100000;
                prev_state = State1_279;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_141)
            begin
                // Must create 281/512*Vdd
                Q = 30'b111100010000000000000000010000;
                prev_state = State1_281;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_141)
            begin
                // Must create 283/512*Vdd
                Q = 30'b111100010000000000000000100000;
                prev_state = State1_283;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_143)
            begin
                // Must create 285/512*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State1_285;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_143)
            begin
                // Must create 287/512*Vdd
                Q = 30'b110000001000000000001100001000;
                prev_state = State1_287;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_145)
            begin
                // Must create 289/512*Vdd
                Q = 30'b101011000000000100000000010000;
                prev_state = State1_289;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_145)
            begin
                // Must create 291/512*Vdd
                Q = 30'b111100001100000000000000000000;
                prev_state = State1_291;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_147)
            begin
                // Must create 293/512*Vdd
                Q = 30'b111000001000000000000000100100;
                prev_state = State1_293;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_147)
            begin
                // Must create 295/512*Vdd
                Q = 30'b111000001000000000000000110000;
                prev_state = State1_295;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_149)
            begin
                // Must create 297/512*Vdd
                Q = 30'b110010000000000000000010110000;
                prev_state = State1_297;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_149)
            begin
                // Must create 299/512*Vdd
                Q = 30'b101000000000000000000011110000;
                prev_state = State1_299;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_151)
            begin
                // Must create 301/512*Vdd
                Q = 30'b111000000000000000000000111000;
                prev_state = State1_301;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_151)
            begin
                // Must create 303/512*Vdd
                Q = 30'b100100010000000000000000111000;
                prev_state = State1_303;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_153)
            begin
                // Must create 305/512*Vdd
                Q = 30'b111000000000000000000000000111;
                prev_state = State1_305;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_153)
            begin
                // Must create 307/512*Vdd
                Q = 30'b100000001100000000000000000111;
                prev_state = State1_307;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_155)
            begin
                // Must create 309/512*Vdd
                Q = 30'b101100000000000000000000000111;
                prev_state = State1_309;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_155)
            begin
                // Must create 311/512*Vdd
                Q = 30'b101100000000000000001000000110;
                prev_state = State1_311;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_157)
            begin
                // Must create 313/512*Vdd
                Q = 30'b100011000000000000100010100000;
                prev_state = State1_313;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_157)
            begin
                // Must create 315/512*Vdd
                Q = 30'b111000000000000000000000111000;
                prev_state = State1_315;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_159)
            begin
                // Must create 317/512*Vdd
                Q = 30'b110010000000000000000000111000;
                prev_state = State1_317;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_159)
            begin
                // Must create 319/512*Vdd
                Q = 30'b100000001000000100000000100110;
                prev_state = State1_319;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_161)
            begin
                // Must create 321/512*Vdd
                Q = 30'b100000000000000000001000000000;
                prev_state = State1_321;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_161)
            begin
                // Must create 323/512*Vdd
                Q = 30'b101000010000000010001000000010;
                prev_state = State1_323;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_163)
            begin
                // Must create 325/512*Vdd
                Q = 30'b111000000000000010000000000011;
                prev_state = State1_325;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_163)
            begin
                // Must create 327/512*Vdd
                Q = 30'b111100000000000010000000000010;
                prev_state = State1_327;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_165)
            begin
                // Must create 329/512*Vdd
                Q = 30'b111101000000000000010000000000;
                prev_state = State1_329;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_165)
            begin
                // Must create 331/512*Vdd
                Q = 30'b111101100000000000000000000000;
                prev_state = State1_331;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_167)
            begin
                // Must create 333/512*Vdd
                Q = 30'b111101100000000000000000000000;
                prev_state = State1_333;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_167)
            begin
                // Must create 335/512*Vdd
                Q = 30'b100101100000000001000000000100;
                prev_state = State1_335;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_169)
            begin
                // Must create 337/512*Vdd
                Q = 30'b110000010000000000010000000011;
                prev_state = State1_337;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_169)
            begin
                // Must create 339/512*Vdd
                Q = 30'b101100010000000000000000000011;
                prev_state = State1_339;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_171)
            begin
                // Must create 341/512*Vdd
                Q = 30'b111000010000000000000000000011;
                prev_state = State1_341;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_171)
            begin
                // Must create 343/512*Vdd
                Q = 30'b111000010000000001000000000010;
                prev_state = State1_343;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_173)
            begin
                // Must create 345/512*Vdd
                Q = 30'b111100000000000000100000000010;
                prev_state = State1_345;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_173)
            begin
                // Must create 347/512*Vdd
                Q = 30'b111000000000000000100000000011;
                prev_state = State1_347;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_175)
            begin
                // Must create 349/512*Vdd
                Q = 30'b101000010000000000100010000010;
                prev_state = State1_349;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_175)
            begin
                // Must create 351/512*Vdd
                Q = 30'b100000000000000000000010000000;
                prev_state = State1_351;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_177)
            begin
                // Must create 353/512*Vdd
                Q = 30'b100000000000000000000010000000;
                prev_state = State1_353;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_177)
            begin
                // Must create 355/512*Vdd
                Q = 30'b111100000000000001100000000000;
                prev_state = State1_355;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_179)
            begin
                // Must create 357/512*Vdd
                Q = 30'b111110000000000000001000000000;
                prev_state = State1_357;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_179)
            begin
                // Must create 359/512*Vdd
                Q = 30'b111110000000000000000000100000;
                prev_state = State1_359;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_181)
            begin
                // Must create 361/512*Vdd
                Q = 30'b111000000000000001110000000000;
                prev_state = State1_361;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_181)
            begin
                // Must create 363/512*Vdd
                Q = 30'b111110000000000100000000000000;
                prev_state = State1_363;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_183)
            begin
                // Must create 365/512*Vdd
                Q = 30'b100100000000000110001000010000;
                prev_state = State1_365;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_183)
            begin
                // Must create 367/512*Vdd
                Q = 30'b100010000000000000000000000000;
                prev_state = State1_367;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_185)
            begin
                // Must create 369/512*Vdd
                Q = 30'b100010000000000000000000000000;
                prev_state = State1_369;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_185)
            begin
                // Must create 371/512*Vdd
                Q = 30'b111100000000000100100000000000;
                prev_state = State1_371;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_187)
            begin
                // Must create 373/512*Vdd
                Q = 30'b111100000000000001010000000000;
                prev_state = State1_373;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_187)
            begin
                // Must create 375/512*Vdd
                Q = 30'b111100000000000001100000000000;
                prev_state = State1_375;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_189)
            begin
                // Must create 377/512*Vdd
                Q = 30'b110000000000000001011100000000;
                prev_state = State1_377;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_189)
            begin
                // Must create 379/512*Vdd
                Q = 30'b100000000000000001011100001000;
                prev_state = State1_379;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_191)
            begin
                // Must create 381/512*Vdd
                Q = 30'b100000000000000101011100000000;
                prev_state = State1_381;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_191)
            begin
                // Must create 383/512*Vdd
                Q = 30'b100000000000000110000000000010;
                prev_state = State1_383;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_193)
            begin
                // Must create 385/512*Vdd
                Q = 30'b100000000000000001000000000000;
                prev_state = State1_385;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_193)
            begin
                // Must create 387/512*Vdd
                Q = 30'b100100000000000111100000000000;
                prev_state = State1_387;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_195)
            begin
                // Must create 389/512*Vdd
                Q = 30'b110100000000000111000000000000;
                prev_state = State1_389;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_195)
            begin
                // Must create 391/512*Vdd
                Q = 30'b110100000000000001000000100100;
                prev_state = State1_391;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_197)
            begin
                // Must create 393/512*Vdd
                Q = 30'b110100000000000001000000001100;
                prev_state = State1_393;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_197)
            begin
                // Must create 395/512*Vdd
                Q = 30'b110100000000000100010000001000;
                prev_state = State1_395;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_199)
            begin
                // Must create 397/512*Vdd
                Q = 30'b111000000000000000010000110000;
                prev_state = State1_397;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_199)
            begin
                // Must create 399/512*Vdd
                Q = 30'b100000000000000000011000110100;
                prev_state = State1_399;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_201)
            begin
                // Must create 401/512*Vdd
                Q = 30'b101000000000000110001000000001;
                prev_state = State1_401;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_201)
            begin
                // Must create 403/512*Vdd
                Q = 30'b110100000000000100010000100000;
                prev_state = State1_403;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_203)
            begin
                // Must create 405/512*Vdd
                Q = 30'b110100000000000100010000100000;
                prev_state = State1_405;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_203)
            begin
                // Must create 407/512*Vdd
                Q = 30'b111100000000000100010000000000;
                prev_state = State1_407;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_205)
            begin
                // Must create 409/512*Vdd
                Q = 30'b111100000000000000000100000010;
                prev_state = State1_409;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_205)
            begin
                // Must create 411/512*Vdd
                Q = 30'b111000000000000101000100000000;
                prev_state = State1_411;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_207)
            begin
                // Must create 413/512*Vdd
                Q = 30'b111000000000000100000011000000;
                prev_state = State1_413;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_207)
            begin
                // Must create 415/512*Vdd
                Q = 30'b100000000000000000000010000000;
                prev_state = State1_415;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_209)
            begin
                // Must create 417/512*Vdd
                Q = 30'b100000000000000000000010000000;
                prev_state = State1_417;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_209)
            begin
                // Must create 419/512*Vdd
                Q = 30'b111000000000000100100100000000;
                prev_state = State1_419;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_211)
            begin
                // Must create 421/512*Vdd
                Q = 30'b111000000000000101001000000000;
                prev_state = State1_421;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_211)
            begin
                // Must create 423/512*Vdd
                Q = 30'b111000000000000101000000100000;
                prev_state = State1_423;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_213)
            begin
                // Must create 425/512*Vdd
                Q = 30'b100000000000000001100001010100;
                prev_state = State1_425;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_213)
            begin
                // Must create 427/512*Vdd
                Q = 30'b110000000000000100011100000000;
                prev_state = State1_427;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_215)
            begin
                // Must create 429/512*Vdd
                Q = 30'b100000000000000101011010000000;
                prev_state = State1_429;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_215)
            begin
                // Must create 431/512*Vdd
                Q = 30'b111000000000000001000000000000;
                prev_state = State1_431;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_217)
            begin
                // Must create 433/512*Vdd
                Q = 30'b100000000000000000001001001110;
                prev_state = State1_433;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_217)
            begin
                // Must create 435/512*Vdd
                Q = 30'b111000000000000000000000001110;
                prev_state = State1_435;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_219)
            begin
                // Must create 437/512*Vdd
                Q = 30'b111000000000000000000000001110;
                prev_state = State1_437;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_219)
            begin
                // Must create 439/512*Vdd
                Q = 30'b111000000000000000010000001100;
                prev_state = State1_439;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_221)
            begin
                // Must create 441/512*Vdd
                Q = 30'b110000000000000000001100000000;
                prev_state = State1_441;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_221)
            begin
                // Must create 443/512*Vdd
                Q = 30'b111000000000000000010011000000;
                prev_state = State1_443;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_223)
            begin
                // Must create 445/512*Vdd
                Q = 30'b111000000000000001000011000000;
                prev_state = State1_445;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_223)
            begin
                // Must create 447/512*Vdd
                Q = 30'b110000000000000000100000000010;
                prev_state = State1_447;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_225)
            begin
                // Must create 449/512*Vdd
                Q = 30'b110000000000000000000000000000;
                prev_state = State1_449;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_225)
            begin
                // Must create 451/512*Vdd
                Q = 30'b010000000000000110100010100000;
                prev_state = State1_451;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_227)
            begin
                // Must create 453/512*Vdd
                Q = 30'b010000000000000101000000111000;
                prev_state = State1_453;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_227)
            begin
                // Must create 455/512*Vdd
                Q = 30'b010000000000000000000100000000;
                prev_state = State1_455;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_229)
            begin
                // Must create 457/512*Vdd
                Q = 30'b110000000000000100010001100000;
                prev_state = State1_457;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_229)
            begin
                // Must create 459/512*Vdd
                Q = 30'b110000000000000101001000100000;
                prev_state = State1_459;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_231)
            begin
                // Must create 461/512*Vdd
                Q = 30'b110000000000000101101000000000;
                prev_state = State1_461;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_231)
            begin
                // Must create 463/512*Vdd
                Q = 30'b110000000000000000000000110000;
                prev_state = State1_463;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_233)
            begin
                // Must create 465/512*Vdd
                Q = 30'b100000000000000001010010000000;
                prev_state = State1_465;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_233)
            begin
                // Must create 467/512*Vdd
                Q = 30'b110000000000000101001001000000;
                prev_state = State1_467;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_235)
            begin
                // Must create 469/512*Vdd
                Q = 30'b110000000000000100001001001000;
                prev_state = State1_469;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_235)
            begin
                // Must create 471/512*Vdd
                Q = 30'b110000000000000100000100001100;
                prev_state = State1_471;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_237)
            begin
                // Must create 473/512*Vdd
                Q = 30'b110000000000000000000000110000;
                prev_state = State1_473;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_237)
            begin
                // Must create 475/512*Vdd
                Q = 30'b110000000000000100001101000000;
                prev_state = State1_475;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_239)
            begin
                // Must create 477/512*Vdd
                Q = 30'b110000000000000100001000110000;
                prev_state = State1_477;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_239)
            begin
                // Must create 479/512*Vdd
                Q = 30'b100000000000000000000100000000;
                prev_state = State1_479;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_241)
            begin
                // Must create 481/512*Vdd
                Q = 30'b100000000000000000000100000000;
                prev_state = State1_481;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_241)
            begin
                // Must create 483/512*Vdd
                Q = 30'b110000000000000001011000100000;
                prev_state = State1_483;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_243)
            begin
                // Must create 485/512*Vdd
                Q = 30'b110000000000000001001101000000;
                prev_state = State1_485;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_243)
            begin
                // Must create 487/512*Vdd
                Q = 30'b110000000000000000000000001100;
                prev_state = State1_487;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_245)
            begin
                // Must create 489/512*Vdd
                Q = 30'b010000000000000001001010000000;
                prev_state = State1_489;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_245)
            begin
                // Must create 491/512*Vdd
                Q = 30'b010000000000000001001100011000;
                prev_state = State1_491;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_247)
            begin
                // Must create 493/512*Vdd
                Q = 30'b010000000000000001000001011100;
                prev_state = State1_493;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_247)
            begin
                // Must create 495/512*Vdd
                Q = 30'b010000000000000000000001000000;
                prev_state = State1_495;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_249)
            begin
                // Must create 497/512*Vdd
                Q = 30'b110000000000000000000000010111;
                prev_state = State1_497;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_249)
            begin
                // Must create 499/512*Vdd
                Q = 30'b010000000000000000001000011000;
                prev_state = State1_499;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_251)
            begin
                // Must create 501/512*Vdd
                Q = 30'b010000000000000000000010011011;
                prev_state = State1_501;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_251)
            begin
                // Must create 503/512*Vdd
                Q = 30'b010000000000000000001100011010;
                prev_state = State1_503;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_253)
            begin
                // Must create 505/512*Vdd
                Q = 30'b010000000000000000001001011010;
                prev_state = State1_505;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_253)
            begin
                // Must create 507/512*Vdd
                Q = 30'b010000000000000000001000010010;
                prev_state = State1_507;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State2_255)
            begin
                // Must create 509/512*Vdd
                Q = 30'b010000000000000000000000010110;
                prev_state = State1_509;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State2_255)
            begin
                // Must create 511/512*Vdd
                Q = 30'b010000000000000000000000000010;
                prev_state = State1_511;
            end
    end
  State0:
    begin
        next_state = INIT;
        data_clk = 1'b1;
        get_comp = 1'b1;
        if (comp_reg == 1'b0 && prev_state_reg == State1_1)
            begin
                // Must create 1/1024*Vdd
                Q = 30'b010000000000001000000000000000;
                prev_state = State0_1;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_1)
            begin
                // Must create 3/1024*Vdd
                Q = 30'b010000000001011000000000000000;
                prev_state = State0_3;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_3)
            begin
                // Must create 5/1024*Vdd
                Q = 30'b010000000011001000000000000000;
                prev_state = State0_5;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_3)
            begin
                // Must create 7/1024*Vdd
                Q = 30'b010000000001000000000000000000;
                prev_state = State0_7;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_5)
            begin
                // Must create 9/1024*Vdd
                Q = 30'b010001000011101000000000000000;
                prev_state = State0_9;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_5)
            begin
                // Must create 11/1024*Vdd
                Q = 30'b010001000001100000000000000000;
                prev_state = State0_11;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_7)
            begin
                // Must create 13/1024*Vdd
                Q = 30'b010000000000100000000000000000;
                prev_state = State0_13;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_7)
            begin
                // Must create 15/1024*Vdd
                Q = 30'b010001000100001000000000000000;
                prev_state = State0_15;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_9)
            begin
                // Must create 17/1024*Vdd
                Q = 30'b010001001000001000000000000000;
                prev_state = State0_17;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_9)
            begin
                // Must create 19/1024*Vdd
                Q = 30'b010000000000100000000000000000;
                prev_state = State0_19;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_11)
            begin
                // Must create 21/1024*Vdd
                Q = 30'b010001110010100000000000000000;
                prev_state = State0_21;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_11)
            begin
                // Must create 23/1024*Vdd
                Q = 30'b010001111010000000000000000000;
                prev_state = State0_23;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_13)
            begin
                // Must create 25/1024*Vdd
                Q = 30'b010000110100110000000000000000;
                prev_state = State0_25;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_13)
            begin
                // Must create 27/1024*Vdd
                Q = 30'b010001101000000000000000000000;
                prev_state = State0_27;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_15)
            begin
                // Must create 29/1024*Vdd
                Q = 30'b110001101010000000000000000000;
                prev_state = State0_29;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_15)
            begin
                // Must create 31/1024*Vdd
                Q = 30'b100000000100000000000000000000;
                prev_state = State0_31;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_17)
            begin
                // Must create 33/1024*Vdd
                Q = 30'b010000000100000000000000000000;
                prev_state = State0_33;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_17)
            begin
                // Must create 35/1024*Vdd
                Q = 30'b011000001100000000000000000000;
                prev_state = State0_35;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_19)
            begin
                // Must create 37/1024*Vdd
                Q = 30'b011000001111000000000000000000;
                prev_state = State0_37;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_19)
            begin
                // Must create 39/1024*Vdd
                Q = 30'b011000001100011000000000000000;
                prev_state = State0_39;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_21)
            begin
                // Must create 41/1024*Vdd
                Q = 30'b011001001000011000000000000000;
                prev_state = State0_41;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_21)
            begin
                // Must create 43/1024*Vdd
                Q = 30'b011001100010010000000000000000;
                prev_state = State0_43;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_23)
            begin
                // Must create 45/1024*Vdd
                Q = 30'b011001100011000000000000000000;
                prev_state = State0_45;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_23)
            begin
                // Must create 47/1024*Vdd
                Q = 30'b010000000000010000000000000000;
                prev_state = State0_47;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_25)
            begin
                // Must create 49/1024*Vdd
                Q = 30'b100000000000010000000000000000;
                prev_state = State0_49;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_25)
            begin
                // Must create 51/1024*Vdd
                Q = 30'b111001001001000000000000000000;
                prev_state = State0_51;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_27)
            begin
                // Must create 53/1024*Vdd
                Q = 30'b111001100001000000000000000000;
                prev_state = State0_53;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_27)
            begin
                // Must create 55/1024*Vdd
                Q = 30'b111000010011000000000000000000;
                prev_state = State0_55;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_29)
            begin
                // Must create 57/1024*Vdd
                Q = 30'b110000001010000000000000000000;
                prev_state = State0_57;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_29)
            begin
                // Must create 59/1024*Vdd
                Q = 30'b111000000001110000000000000000;
                prev_state = State0_59;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_31)
            begin
                // Must create 61/1024*Vdd
                Q = 30'b100010010101100000000000000000;
                prev_state = State0_61;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_31)
            begin
                // Must create 63/1024*Vdd
                Q = 30'b100000010000000000000000000000;
                prev_state = State0_63;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_33)
            begin
                // Must create 65/1024*Vdd
                Q = 30'b100000010000000000000000000000;
                prev_state = State0_65;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_33)
            begin
                // Must create 67/1024*Vdd
                Q = 30'b100000010011101000000000000000;
                prev_state = State0_67;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_35)
            begin
                // Must create 69/1024*Vdd
                Q = 30'b110001000000101100000000000000;
                prev_state = State0_69;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_35)
            begin
                // Must create 71/1024*Vdd
                Q = 30'b110000000100010000000000000000;
                prev_state = State0_71;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_37)
            begin
                // Must create 73/1024*Vdd
                Q = 30'b110001010010010000000000000000;
                prev_state = State0_73;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_37)
            begin
                // Must create 75/1024*Vdd
                Q = 30'b110001101010000000000000000000;
                prev_state = State0_75;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_39)
            begin
                // Must create 77/1024*Vdd
                Q = 30'b110001001110000000000000000000;
                prev_state = State0_77;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_39)
            begin
                // Must create 79/1024*Vdd
                Q = 30'b100000000000100000000000000000;
                prev_state = State0_79;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_41)
            begin
                // Must create 81/1024*Vdd
                Q = 30'b100000011111000000000000000000;
                prev_state = State0_81;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_41)
            begin
                // Must create 83/1024*Vdd
                Q = 30'b110001001110000000000000000000;
                prev_state = State0_83;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_43)
            begin
                // Must create 85/1024*Vdd
                Q = 30'b110001001100100000000000000000;
                prev_state = State0_85;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_43)
            begin
                // Must create 87/1024*Vdd
                Q = 30'b100000000001000000000000000000;
                prev_state = State0_87;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_45)
            begin
                // Must create 89/1024*Vdd
                Q = 30'b110000000011000000000000000000;
                prev_state = State0_89;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_45)
            begin
                // Must create 91/1024*Vdd
                Q = 30'b111000100000110000000000000000;
                prev_state = State0_91;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_47)
            begin
                // Must create 93/1024*Vdd
                Q = 30'b101011100000100000000000000000;
                prev_state = State0_93;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_47)
            begin
                // Must create 95/1024*Vdd
                Q = 30'b100000000000000100000000000000;
                prev_state = State0_95;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_49)
            begin
                // Must create 97/1024*Vdd
                Q = 30'b100000000000000100000000000000;
                prev_state = State0_97;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_49)
            begin
                // Must create 99/1024*Vdd
                Q = 30'b110100000110100000000000000000;
                prev_state = State0_99;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_51)
            begin
                // Must create 101/1024*Vdd
                Q = 30'b111000000100110000000000000000;
                prev_state = State0_101;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_51)
            begin
                // Must create 103/1024*Vdd
                Q = 30'b100010000111000100000000000000;
                prev_state = State0_103;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_53)
            begin
                // Must create 105/1024*Vdd
                Q = 30'b111000001101000000000000000000;
                prev_state = State0_105;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_53)
            begin
                // Must create 107/1024*Vdd
                Q = 30'b111001100100000000000000000000;
                prev_state = State0_107;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_55)
            begin
                // Must create 109/1024*Vdd
                Q = 30'b111001110000000000000000000000;
                prev_state = State0_109;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_55)
            begin
                // Must create 111/1024*Vdd
                Q = 30'b100101000001100100000000000000;
                prev_state = State0_111;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_57)
            begin
                // Must create 113/1024*Vdd
                Q = 30'b010000000100000000000000000000;
                prev_state = State0_113;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_57)
            begin
                // Must create 115/1024*Vdd
                Q = 30'b011101100100000000000000000000;
                prev_state = State0_115;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_59)
            begin
                // Must create 117/1024*Vdd
                Q = 30'b011101110000000000000000000000;
                prev_state = State0_117;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_59)
            begin
                // Must create 119/1024*Vdd
                Q = 30'b111101100000000000000000000000;
                prev_state = State0_119;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_61)
            begin
                // Must create 121/1024*Vdd
                Q = 30'b011101000000011000000000000000;
                prev_state = State0_121;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_61)
            begin
                // Must create 123/1024*Vdd
                Q = 30'b011100000000011010000000000000;
                prev_state = State0_123;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_63)
            begin
                // Must create 125/1024*Vdd
                Q = 30'b101010000000111000000000000000;
                prev_state = State0_125;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_63)
            begin
                // Must create 127/1024*Vdd
                Q = 30'b100010000000000000000000000000;
                prev_state = State0_127;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_65)
            begin
                // Must create 129/1024*Vdd
                Q = 30'b100010000000000000000000000000;
                prev_state = State0_129;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_65)
            begin
                // Must create 131/1024*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State0_131;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_67)
            begin
                // Must create 133/1024*Vdd
                Q = 30'b111011001000000000000000000000;
                prev_state = State0_133;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_67)
            begin
                // Must create 135/1024*Vdd
                Q = 30'b111010100000000001000000000000;
                prev_state = State0_135;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_69)
            begin
                // Must create 137/1024*Vdd
                Q = 30'b101000110001100000000000000000;
                prev_state = State0_137;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_69)
            begin
                // Must create 139/1024*Vdd
                Q = 30'b110011101000000000000000000000;
                prev_state = State0_139;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_71)
            begin
                // Must create 141/1024*Vdd
                Q = 30'b110001101100000000000000000000;
                prev_state = State0_141;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_71)
            begin
                // Must create 143/1024*Vdd
                Q = 30'b100000000010000000000000000000;
                prev_state = State0_143;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_73)
            begin
                // Must create 145/1024*Vdd
                Q = 30'b110000010010000000000000000000;
                prev_state = State0_145;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_73)
            begin
                // Must create 147/1024*Vdd
                Q = 30'b111001100001000000000000000000;
                prev_state = State0_147;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_75)
            begin
                // Must create 149/1024*Vdd
                Q = 30'b111001100001000000000000000000;
                prev_state = State0_149;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_75)
            begin
                // Must create 151/1024*Vdd
                Q = 30'b111001100100000000000000000000;
                prev_state = State0_151;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_77)
            begin
                // Must create 153/1024*Vdd
                Q = 30'b111001101000000000000000000000;
                prev_state = State0_153;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_77)
            begin
                // Must create 155/1024*Vdd
                Q = 30'b111001001001000000000000000000;
                prev_state = State0_155;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_79)
            begin
                // Must create 157/1024*Vdd
                Q = 30'b111001100000100000000000000000;
                prev_state = State0_157;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_79)
            begin
                // Must create 159/1024*Vdd
                Q = 30'b100000000100000000000000000000;
                prev_state = State0_159;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_81)
            begin
                // Must create 161/1024*Vdd
                Q = 30'b100000000100000000000000000000;
                prev_state = State0_161;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_81)
            begin
                // Must create 163/1024*Vdd
                Q = 30'b111000001000100100000000000000;
                prev_state = State0_163;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_83)
            begin
                // Must create 165/1024*Vdd
                Q = 30'b101010000000100101000000000000;
                prev_state = State0_165;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_83)
            begin
                // Must create 167/1024*Vdd
                Q = 30'b110000000000111010000000000000;
                prev_state = State0_167;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_85)
            begin
                // Must create 169/1024*Vdd
                Q = 30'b110011000001000100000000000000;
                prev_state = State0_169;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_85)
            begin
                // Must create 171/1024*Vdd
                Q = 30'b110010110000000100000000000000;
                prev_state = State0_171;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_87)
            begin
                // Must create 173/1024*Vdd
                Q = 30'b101110110000000000000000000000;
                prev_state = State0_173;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_87)
            begin
                // Must create 175/1024*Vdd
                Q = 30'b100000000000000100000000000000;
                prev_state = State0_175;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_89)
            begin
                // Must create 177/1024*Vdd
                Q = 30'b100000001010110010000000000000;
                prev_state = State0_177;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_89)
            begin
                // Must create 179/1024*Vdd
                Q = 30'b111000000011000100000000000000;
                prev_state = State0_179;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_91)
            begin
                // Must create 181/1024*Vdd
                Q = 30'b111000000011000100000000000000;
                prev_state = State0_181;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_91)
            begin
                // Must create 183/1024*Vdd
                Q = 30'b111000001011000000000000000000;
                prev_state = State0_183;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_93)
            begin
                // Must create 185/1024*Vdd
                Q = 30'b110000110000000000000000000000;
                prev_state = State0_185;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_93)
            begin
                // Must create 187/1024*Vdd
                Q = 30'b111000000011000100000000000000;
                prev_state = State0_187;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_95)
            begin
                // Must create 189/1024*Vdd
                Q = 30'b100100000111000001000000000000;
                prev_state = State0_189;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_95)
            begin
                // Must create 191/1024*Vdd
                Q = 30'b100000000000000001000000000000;
                prev_state = State0_191;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_97)
            begin
                // Must create 193/1024*Vdd
                Q = 30'b100000000000000001000000000000;
                prev_state = State0_193;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_97)
            begin
                // Must create 195/1024*Vdd
                Q = 30'b110000001000000001000000000000;
                prev_state = State0_195;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_99)
            begin
                // Must create 197/1024*Vdd
                Q = 30'b100000010000000000000000000000;
                prev_state = State0_197;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_99)
            begin
                // Must create 199/1024*Vdd
                Q = 30'b100000100000000000000000000000;
                prev_state = State0_199;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_101)
            begin
                // Must create 201/1024*Vdd
                Q = 30'b111000101000000100000000000000;
                prev_state = State0_201;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_101)
            begin
                // Must create 203/1024*Vdd
                Q = 30'b111001010000000100000000000000;
                prev_state = State0_203;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_103)
            begin
                // Must create 205/1024*Vdd
                Q = 30'b111001000000110000000000000000;
                prev_state = State0_205;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_103)
            begin
                // Must create 207/1024*Vdd
                Q = 30'b100001100100110000000000000000;
                prev_state = State0_207;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_105)
            begin
                // Must create 209/1024*Vdd
                Q = 30'b100000100010110100000000000000;
                prev_state = State0_209;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_105)
            begin
                // Must create 211/1024*Vdd
                Q = 30'b111000000000110100000000000000;
                prev_state = State0_211;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_107)
            begin
                // Must create 213/1024*Vdd
                Q = 30'b111000000000110100000000000000;
                prev_state = State0_213;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_107)
            begin
                // Must create 215/1024*Vdd
                Q = 30'b111000000001110000000000000000;
                prev_state = State0_215;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_109)
            begin
                // Must create 217/1024*Vdd
                Q = 30'b111100000000100100000000000000;
                prev_state = State0_217;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_109)
            begin
                // Must create 219/1024*Vdd
                Q = 30'b111100000000110000000000000000;
                prev_state = State0_219;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_111)
            begin
                // Must create 221/1024*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State0_221;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_111)
            begin
                // Must create 223/1024*Vdd
                Q = 30'b100010000001000000100000000000;
                prev_state = State0_223;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_113)
            begin
                // Must create 225/1024*Vdd
                Q = 30'b111100011000000000000000000000;
                prev_state = State0_225;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_113)
            begin
                // Must create 227/1024*Vdd
                Q = 30'b110011100010000000000000000000;
                prev_state = State0_227;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_115)
            begin
                // Must create 229/1024*Vdd
                Q = 30'b110011000100000000100000000000;
                prev_state = State0_229;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_115)
            begin
                // Must create 231/1024*Vdd
                Q = 30'b110011000100000100000000000000;
                prev_state = State0_231;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_117)
            begin
                // Must create 233/1024*Vdd
                Q = 30'b100000000000100000000000000000;
                prev_state = State0_233;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_117)
            begin
                // Must create 235/1024*Vdd
                Q = 30'b110010000110000100000000000000;
                prev_state = State0_235;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_119)
            begin
                // Must create 237/1024*Vdd
                Q = 30'b111000000111000000000000000000;
                prev_state = State0_237;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_119)
            begin
                // Must create 239/1024*Vdd
                Q = 30'b100100000111100000000000000000;
                prev_state = State0_239;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_121)
            begin
                // Must create 241/1024*Vdd
                Q = 30'b100000000101110010000000000000;
                prev_state = State0_241;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_121)
            begin
                // Must create 243/1024*Vdd
                Q = 30'b111000000100110000000000000000;
                prev_state = State0_243;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_123)
            begin
                // Must create 245/1024*Vdd
                Q = 30'b111010000100000100000000000000;
                prev_state = State0_245;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_123)
            begin
                // Must create 247/1024*Vdd
                Q = 30'b111100000000000110000000000000;
                prev_state = State0_247;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_125)
            begin
                // Must create 249/1024*Vdd
                Q = 30'b100000000000000010000000000000;
                prev_state = State0_249;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_125)
            begin
                // Must create 251/1024*Vdd
                Q = 30'b110000000000000000000000000000;
                prev_state = State0_251;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_127)
            begin
                // Must create 253/1024*Vdd
                Q = 30'b101110000000000000000000000000;
                prev_state = State0_253;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_127)
            begin
                // Must create 255/1024*Vdd
                Q = 30'b100100000000000000000000000000;
                prev_state = State0_255;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_129)
            begin
                // Must create 257/1024*Vdd
                Q = 30'b100100000000000000000000000000;
                prev_state = State0_257;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_129)
            begin
                // Must create 259/1024*Vdd
                Q = 30'b100100110000110000000000000000;
                prev_state = State0_259;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_131)
            begin
                // Must create 261/1024*Vdd
                Q = 30'b100100110001100000000000000000;
                prev_state = State0_261;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_131)
            begin
                // Must create 263/1024*Vdd
                Q = 30'b100100111000000000100000000000;
                prev_state = State0_263;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_133)
            begin
                // Must create 265/1024*Vdd
                Q = 30'b100100111010000000000000000000;
                prev_state = State0_265;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_133)
            begin
                // Must create 267/1024*Vdd
                Q = 30'b100000111010000000010000000000;
                prev_state = State0_267;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_135)
            begin
                // Must create 269/1024*Vdd
                Q = 30'b110000101010000000010000000000;
                prev_state = State0_269;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_135)
            begin
                // Must create 271/1024*Vdd
                Q = 30'b101000001010000000110000000000;
                prev_state = State0_271;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_137)
            begin
                // Must create 273/1024*Vdd
                Q = 30'b100001001101000100000000000000;
                prev_state = State0_273;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_137)
            begin
                // Must create 275/1024*Vdd
                Q = 30'b111000001010000000010000000000;
                prev_state = State0_275;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_139)
            begin
                // Must create 277/1024*Vdd
                Q = 30'b111000001010000000010000000000;
                prev_state = State0_277;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_139)
            begin
                // Must create 279/1024*Vdd
                Q = 30'b111001001010000000000000000000;
                prev_state = State0_279;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_141)
            begin
                // Must create 281/1024*Vdd
                Q = 30'b111000000011000100000000000000;
                prev_state = State0_281;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_141)
            begin
                // Must create 283/1024*Vdd
                Q = 30'b111000000001000101000000000000;
                prev_state = State0_283;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_143)
            begin
                // Must create 285/1024*Vdd
                Q = 30'b100100001101000100000000000000;
                prev_state = State0_285;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_143)
            begin
                // Must create 287/1024*Vdd
                Q = 30'b100000000100000000000000000000;
                prev_state = State0_287;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_145)
            begin
                // Must create 289/1024*Vdd
                Q = 30'b100000000100000000000000000000;
                prev_state = State0_289;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_145)
            begin
                // Must create 291/1024*Vdd
                Q = 30'b100010001101000010000000000000;
                prev_state = State0_291;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_147)
            begin
                // Must create 293/1024*Vdd
                Q = 30'b100010001001000010010000000000;
                prev_state = State0_293;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_147)
            begin
                // Must create 295/1024*Vdd
                Q = 30'b110010001001000010000000000000;
                prev_state = State0_295;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_149)
            begin
                // Must create 297/1024*Vdd
                Q = 30'b111100000100000001000000000000;
                prev_state = State0_297;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_149)
            begin
                // Must create 299/1024*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State0_299;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_151)
            begin
                // Must create 301/1024*Vdd
                Q = 30'b111010000010000100000000000000;
                prev_state = State0_301;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_151)
            begin
                // Must create 303/1024*Vdd
                Q = 30'b100010001010000101000000000000;
                prev_state = State0_303;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_153)
            begin
                // Must create 305/1024*Vdd
                Q = 30'b100100001010000100100000000000;
                prev_state = State0_305;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_153)
            begin
                // Must create 307/1024*Vdd
                Q = 30'b111100110000000000000000000000;
                prev_state = State0_307;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_155)
            begin
                // Must create 309/1024*Vdd
                Q = 30'b111100110000000000000000000000;
                prev_state = State0_309;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_155)
            begin
                // Must create 311/1024*Vdd
                Q = 30'b111100101000000000000000000000;
                prev_state = State0_311;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_157)
            begin
                // Must create 313/1024*Vdd
                Q = 30'b110001000000000001000000000000;
                prev_state = State0_313;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_157)
            begin
                // Must create 315/1024*Vdd
                Q = 30'b111000010100000000100000000000;
                prev_state = State0_315;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_159)
            begin
                // Must create 317/1024*Vdd
                Q = 30'b100100110100000000010000000000;
                prev_state = State0_317;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_159)
            begin
                // Must create 319/1024*Vdd
                Q = 30'b100000000000000000010000000000;
                prev_state = State0_319;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_161)
            begin
                // Must create 321/1024*Vdd
                Q = 30'b100000000000000000010000000000;
                prev_state = State0_321;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_161)
            begin
                // Must create 323/1024*Vdd
                Q = 30'b100100001000000000010000000000;
                prev_state = State0_323;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_163)
            begin
                // Must create 325/1024*Vdd
                Q = 30'b100110001000010000010000000000;
                prev_state = State0_325;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_163)
            begin
                // Must create 327/1024*Vdd
                Q = 30'b110110000000000000010010000000;
                prev_state = State0_327;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_165)
            begin
                // Must create 329/1024*Vdd
                Q = 30'b111110010000000000000000000000;
                prev_state = State0_329;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_165)
            begin
                // Must create 331/1024*Vdd
                Q = 30'b111110000001000000000000000000;
                prev_state = State0_331;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_167)
            begin
                // Must create 333/1024*Vdd
                Q = 30'b111110000001000000000000000000;
                prev_state = State0_333;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_167)
            begin
                // Must create 335/1024*Vdd
                Q = 30'b100110000101000000000010000000;
                prev_state = State0_335;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_169)
            begin
                // Must create 337/1024*Vdd
                Q = 30'b100011001001000000000010000000;
                prev_state = State0_337;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_169)
            begin
                // Must create 339/1024*Vdd
                Q = 30'b111011000001000000000000000000;
                prev_state = State0_339;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_171)
            begin
                // Must create 341/1024*Vdd
                Q = 30'b111011000001000000000000000000;
                prev_state = State0_341;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_171)
            begin
                // Must create 343/1024*Vdd
                Q = 30'b111011000100000000000000000000;
                prev_state = State0_343;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_173)
            begin
                // Must create 345/1024*Vdd
                Q = 30'b110011000110000000000000000000;
                prev_state = State0_345;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_173)
            begin
                // Must create 347/1024*Vdd
                Q = 30'b100011000110000000001000000000;
                prev_state = State0_347;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_175)
            begin
                // Must create 349/1024*Vdd
                Q = 30'b110011100100000000000000000000;
                prev_state = State0_349;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_175)
            begin
                // Must create 351/1024*Vdd
                Q = 30'b111000100001000001000000000000;
                prev_state = State0_351;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_177)
            begin
                // Must create 353/1024*Vdd
                Q = 30'b110000100000011000000010000000;
                prev_state = State0_353;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_177)
            begin
                // Must create 355/1024*Vdd
                Q = 30'b111011010000000000000000000000;
                prev_state = State0_355;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_179)
            begin
                // Must create 357/1024*Vdd
                Q = 30'b111010000000100100000000000000;
                prev_state = State0_357;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_179)
            begin
                // Must create 359/1024*Vdd
                Q = 30'b111010000000100000000100000000;
                prev_state = State0_359;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_181)
            begin
                // Must create 361/1024*Vdd
                Q = 30'b110010000010100100000000000000;
                prev_state = State0_361;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_181)
            begin
                // Must create 363/1024*Vdd
                Q = 30'b110010000000100100000100000000;
                prev_state = State0_363;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_183)
            begin
                // Must create 365/1024*Vdd
                Q = 30'b110010000000100100000100000000;
                prev_state = State0_365;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_183)
            begin
                // Must create 367/1024*Vdd
                Q = 30'b100000000001100101000100000000;
                prev_state = State0_367;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_185)
            begin
                // Must create 369/1024*Vdd
                Q = 30'b100000000101110000000010000000;
                prev_state = State0_369;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_185)
            begin
                // Must create 371/1024*Vdd
                Q = 30'b110010000001110000000000000000;
                prev_state = State0_371;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_187)
            begin
                // Must create 373/1024*Vdd
                Q = 30'b110010000001110000000000000000;
                prev_state = State0_373;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_187)
            begin
                // Must create 375/1024*Vdd
                Q = 30'b110010100001100000000000000000;
                prev_state = State0_375;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_189)
            begin
                // Must create 377/1024*Vdd
                Q = 30'b110010000000010000100010000000;
                prev_state = State0_377;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_189)
            begin
                // Must create 379/1024*Vdd
                Q = 30'b100010000000011010100000000000;
                prev_state = State0_379;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_191)
            begin
                // Must create 381/1024*Vdd
                Q = 30'b100010000000000001100000000000;
                prev_state = State0_381;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_191)
            begin
                // Must create 383/1024*Vdd
                Q = 30'b100000000000000000100000000000;
                prev_state = State0_383;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_193)
            begin
                // Must create 385/1024*Vdd
                Q = 30'b100000000001000001100000000000;
                prev_state = State0_385;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_193)
            begin
                // Must create 387/1024*Vdd
                Q = 30'b111100000001100000000000000000;
                prev_state = State0_387;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_195)
            begin
                // Must create 389/1024*Vdd
                Q = 30'b111100011000000000000000000000;
                prev_state = State0_389;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_195)
            begin
                // Must create 391/1024*Vdd
                Q = 30'b111110010000000000000000000000;
                prev_state = State0_391;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_197)
            begin
                // Must create 393/1024*Vdd
                Q = 30'b111011000000000001000000000000;
                prev_state = State0_393;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_197)
            begin
                // Must create 395/1024*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State0_395;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_199)
            begin
                // Must create 397/1024*Vdd
                Q = 30'b111110010000000000000000000000;
                prev_state = State0_397;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_199)
            begin
                // Must create 399/1024*Vdd
                Q = 30'b100100000110000000000000000000;
                prev_state = State0_399;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_201)
            begin
                // Must create 401/1024*Vdd
                Q = 30'b100000100000110000100000100000;
                prev_state = State0_401;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_201)
            begin
                // Must create 403/1024*Vdd
                Q = 30'b100011100000110000000000000000;
                prev_state = State0_403;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_203)
            begin
                // Must create 405/1024*Vdd
                Q = 30'b100011100000110000000000000000;
                prev_state = State0_405;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_203)
            begin
                // Must create 407/1024*Vdd
                Q = 30'b100011100001100000000000000000;
                prev_state = State0_407;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_205)
            begin
                // Must create 409/1024*Vdd
                Q = 30'b100010000001110000000100000000;
                prev_state = State0_409;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_205)
            begin
                // Must create 411/1024*Vdd
                Q = 30'b100000000001110000000110000000;
                prev_state = State0_411;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_207)
            begin
                // Must create 413/1024*Vdd
                Q = 30'b110010000001110000000000000000;
                prev_state = State0_413;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_207)
            begin
                // Must create 415/1024*Vdd
                Q = 30'b110011110000000000000000000000;
                prev_state = State0_415;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_209)
            begin
                // Must create 417/1024*Vdd
                Q = 30'b110000100000000001011000000000;
                prev_state = State0_417;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_209)
            begin
                // Must create 419/1024*Vdd
                Q = 30'b110011010010000000000000000000;
                prev_state = State0_419;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_211)
            begin
                // Must create 421/1024*Vdd
                Q = 30'b110010011100000000000000000000;
                prev_state = State0_421;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_211)
            begin
                // Must create 423/1024*Vdd
                Q = 30'b110010011010000000000000000000;
                prev_state = State0_423;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_213)
            begin
                // Must create 425/1024*Vdd
                Q = 30'b100000000000000000000010000000;
                prev_state = State0_425;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_213)
            begin
                // Must create 427/1024*Vdd
                Q = 30'b110010011001000000000000000000;
                prev_state = State0_427;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_215)
            begin
                // Must create 429/1024*Vdd
                Q = 30'b110000011110000000000000000000;
                prev_state = State0_429;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_215)
            begin
                // Must create 431/1024*Vdd
                Q = 30'b100000001110000000001010000000;
                prev_state = State0_431;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_217)
            begin
                // Must create 433/1024*Vdd
                Q = 30'b100001011000000000000011000000;
                prev_state = State0_433;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_217)
            begin
                // Must create 435/1024*Vdd
                Q = 30'b110011011000000000000000000000;
                prev_state = State0_435;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_219)
            begin
                // Must create 437/1024*Vdd
                Q = 30'b110011011000000000000000000000;
                prev_state = State0_437;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_219)
            begin
                // Must create 439/1024*Vdd
                Q = 30'b110011010000000000010000000000;
                prev_state = State0_439;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_221)
            begin
                // Must create 441/1024*Vdd
                Q = 30'b110010010000010001000000000000;
                prev_state = State0_441;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_221)
            begin
                // Must create 443/1024*Vdd
                Q = 30'b110010000000010001000000100000;
                prev_state = State0_443;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_223)
            begin
                // Must create 445/1024*Vdd
                Q = 30'b110010110000010000000000000000;
                prev_state = State0_445;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_223)
            begin
                // Must create 447/1024*Vdd
                Q = 30'b110000000110000010000010000000;
                prev_state = State0_447;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_225)
            begin
                // Must create 449/1024*Vdd
                Q = 30'b101000100000100100000000100000;
                prev_state = State0_449;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_225)
            begin
                // Must create 451/1024*Vdd
                Q = 30'b110000111001000000000000000000;
                prev_state = State0_451;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_227)
            begin
                // Must create 453/1024*Vdd
                Q = 30'b110010001100000000000010000000;
                prev_state = State0_453;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_227)
            begin
                // Must create 455/1024*Vdd
                Q = 30'b110000000010000000000100000000;
                prev_state = State0_455;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_229)
            begin
                // Must create 457/1024*Vdd
                Q = 30'b110010011000000000010000000000;
                prev_state = State0_457;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_229)
            begin
                // Must create 459/1024*Vdd
                Q = 30'b110010011100000000000000000000;
                prev_state = State0_459;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_231)
            begin
                // Must create 461/1024*Vdd
                Q = 30'b110010011100000000000000000000;
                prev_state = State0_461;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_231)
            begin
                // Must create 463/1024*Vdd
                Q = 30'b100000110001000000010001000000;
                prev_state = State0_463;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_233)
            begin
                // Must create 465/1024*Vdd
                Q = 30'b100000011100000000001010000000;
                prev_state = State0_465;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_233)
            begin
                // Must create 467/1024*Vdd
                Q = 30'b110010011100000000000000000000;
                prev_state = State0_467;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_235)
            begin
                // Must create 469/1024*Vdd
                Q = 30'b110011010010000000000000000000;
                prev_state = State0_469;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_235)
            begin
                // Must create 471/1024*Vdd
                Q = 30'b100000000000000000000010000000;
                prev_state = State0_471;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_237)
            begin
                // Must create 473/1024*Vdd
                Q = 30'b110010001000000000011000000000;
                prev_state = State0_473;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_237)
            begin
                // Must create 475/1024*Vdd
                Q = 30'b110010000000000000011001000000;
                prev_state = State0_475;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_239)
            begin
                // Must create 477/1024*Vdd
                Q = 30'b111000010001000000010000000000;
                prev_state = State0_477;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_239)
            begin
                // Must create 479/1024*Vdd
                Q = 30'b100010011010000100000000000000;
                prev_state = State0_479;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_241)
            begin
                // Must create 481/1024*Vdd
                Q = 30'b110000000000010000011000010000;
                prev_state = State0_481;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_241)
            begin
                // Must create 483/1024*Vdd
                Q = 30'b110010011100000000000000000000;
                prev_state = State0_483;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_243)
            begin
                // Must create 485/1024*Vdd
                Q = 30'b110010010000100000000001000000;
                prev_state = State0_485;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_243)
            begin
                // Must create 487/1024*Vdd
                Q = 30'b110010010000100000000000100000;
                prev_state = State0_487;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_245)
            begin
                // Must create 489/1024*Vdd
                Q = 30'b110010000000100000000101000000;
                prev_state = State0_489;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_245)
            begin
                // Must create 491/1024*Vdd
                Q = 30'b110010000000100000000001100000;
                prev_state = State0_491;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_247)
            begin
                // Must create 493/1024*Vdd
                Q = 30'b110010000100110000000000000000;
                prev_state = State0_493;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_247)
            begin
                // Must create 495/1024*Vdd
                Q = 30'b111100010000000000000000001000;
                prev_state = State0_495;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_249)
            begin
                // Must create 497/1024*Vdd
                Q = 30'b100000000011110000000000001000;
                prev_state = State0_497;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_249)
            begin
                // Must create 499/1024*Vdd
                Q = 30'b110010000001110000000000000000;
                prev_state = State0_499;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_251)
            begin
                // Must create 501/1024*Vdd
                Q = 30'b110010000001110000000000000000;
                prev_state = State0_501;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_251)
            begin
                // Must create 503/1024*Vdd
                Q = 30'b101100000101000000000000000100;
                prev_state = State0_503;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_253)
            begin
                // Must create 505/1024*Vdd
                Q = 30'b111001100001000000000000000000;
                prev_state = State0_505;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_253)
            begin
                // Must create 507/1024*Vdd
                Q = 30'b111001100000000000000000000100;
                prev_state = State0_507;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_255)
            begin
                // Must create 509/1024*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State0_509;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_255)
            begin
                // Must create 511/1024*Vdd
                Q = 30'b100100000000000110000000000000;
                prev_state = State0_511;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_257)
            begin
                // Must create 513/1024*Vdd
                Q = 30'b101000000000000110000000000000;
                prev_state = State0_513;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_257)
            begin
                // Must create 515/1024*Vdd
                Q = 30'b111100000000110000000000000000;
                prev_state = State0_515;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_259)
            begin
                // Must create 517/1024*Vdd
                Q = 30'b111000000000100001010000000000;
                prev_state = State0_517;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_259)
            begin
                // Must create 519/1024*Vdd
                Q = 30'b111000001000100001000000000000;
                prev_state = State0_519;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_261)
            begin
                // Must create 521/1024*Vdd
                Q = 30'b100000101000100001100000000000;
                prev_state = State0_521;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_261)
            begin
                // Must create 523/1024*Vdd
                Q = 30'b111000001110000000000000000000;
                prev_state = State0_523;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_263)
            begin
                // Must create 525/1024*Vdd
                Q = 30'b111000001110000000000000000000;
                prev_state = State0_525;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_263)
            begin
                // Must create 527/1024*Vdd
                Q = 30'b100000011110000000000000000001;
                prev_state = State0_527;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_265)
            begin
                // Must create 529/1024*Vdd
                Q = 30'b110010000001000001100000000000;
                prev_state = State0_529;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_265)
            begin
                // Must create 531/1024*Vdd
                Q = 30'b111000100110000000000000000000;
                prev_state = State0_531;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_267)
            begin
                // Must create 533/1024*Vdd
                Q = 30'b111000000100000000000000001100;
                prev_state = State0_533;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_267)
            begin
                // Must create 535/1024*Vdd
                Q = 30'b111000000100000000000000101000;
                prev_state = State0_535;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_269)
            begin
                // Must create 537/1024*Vdd
                Q = 30'b111010000100000000000000000100;
                prev_state = State0_537;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_269)
            begin
                // Must create 539/1024*Vdd
                Q = 30'b111010000100000000000000001000;
                prev_state = State0_539;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_271)
            begin
                // Must create 541/1024*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State0_541;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_271)
            begin
                // Must create 543/1024*Vdd
                Q = 30'b110000000010000000000011000010;
                prev_state = State0_543;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_273)
            begin
                // Must create 545/1024*Vdd
                Q = 30'b101011010000000100000000000000;
                prev_state = State0_545;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_273)
            begin
                // Must create 547/1024*Vdd
                Q = 30'b110110001000000000000010000000;
                prev_state = State0_547;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_275)
            begin
                // Must create 549/1024*Vdd
                Q = 30'b111000000000000000000011001000;
                prev_state = State0_549;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_275)
            begin
                // Must create 551/1024*Vdd
                Q = 30'b111001000000000000000011000000;
                prev_state = State0_551;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_277)
            begin
                // Must create 553/1024*Vdd
                Q = 30'b100000000000000000000000010000;
                prev_state = State0_553;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_277)
            begin
                // Must create 555/1024*Vdd
                Q = 30'b111110010000000000000000000000;
                prev_state = State0_555;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_279)
            begin
                // Must create 557/1024*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State0_557;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_279)
            begin
                // Must create 559/1024*Vdd
                Q = 30'b100011100000000000000001010000;
                prev_state = State0_559;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_281)
            begin
                // Must create 561/1024*Vdd
                Q = 30'b100010001000000000010010001000;
                prev_state = State0_561;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_281)
            begin
                // Must create 563/1024*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State0_563;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_283)
            begin
                // Must create 565/1024*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State0_565;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_283)
            begin
                // Must create 567/1024*Vdd
                Q = 30'b111011000000000000000010000000;
                prev_state = State0_567;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_285)
            begin
                // Must create 569/1024*Vdd
                Q = 30'b110000010000000000000000100000;
                prev_state = State0_569;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_285)
            begin
                // Must create 571/1024*Vdd
                Q = 30'b111000100000000000010000010000;
                prev_state = State0_571;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_287)
            begin
                // Must create 573/1024*Vdd
                Q = 30'b110011101000000000000000000000;
                prev_state = State0_573;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_287)
            begin
                // Must create 575/1024*Vdd
                Q = 30'b100010000100000101000000000100;
                prev_state = State0_575;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_289)
            begin
                // Must create 577/1024*Vdd
                Q = 30'b110000110000000010000000001000;
                prev_state = State0_577;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_289)
            begin
                // Must create 579/1024*Vdd
                Q = 30'b111010000100000000010000000000;
                prev_state = State0_579;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_291)
            begin
                // Must create 581/1024*Vdd
                Q = 30'b111000000000000000011000000010;
                prev_state = State0_581;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_291)
            begin
                // Must create 583/1024*Vdd
                Q = 30'b111010000000000000011000000000;
                prev_state = State0_583;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_293)
            begin
                // Must create 585/1024*Vdd
                Q = 30'b111110000000000000000010000000;
                prev_state = State0_585;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_293)
            begin
                // Must create 587/1024*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State0_587;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_295)
            begin
                // Must create 589/1024*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State0_589;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_295)
            begin
                // Must create 591/1024*Vdd
                Q = 30'b100111000000000000000000001100;
                prev_state = State0_591;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_297)
            begin
                // Must create 593/1024*Vdd
                Q = 30'b100001110000000000000001001000;
                prev_state = State0_593;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_297)
            begin
                // Must create 595/1024*Vdd
                Q = 30'b110011110000000000000000000000;
                prev_state = State0_595;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_299)
            begin
                // Must create 597/1024*Vdd
                Q = 30'b111011000000000000000010000000;
                prev_state = State0_597;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_299)
            begin
                // Must create 599/1024*Vdd
                Q = 30'b100000000000000000000000001000;
                prev_state = State0_599;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_301)
            begin
                // Must create 601/1024*Vdd
                Q = 30'b111011010000000000000000000000;
                prev_state = State0_601;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_301)
            begin
                // Must create 603/1024*Vdd
                Q = 30'b111011100000000000000000000000;
                prev_state = State0_603;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_303)
            begin
                // Must create 605/1024*Vdd
                Q = 30'b111110010000000000000000000000;
                prev_state = State0_605;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_303)
            begin
                // Must create 607/1024*Vdd
                Q = 30'b110000000000000000011011000000;
                prev_state = State0_607;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_305)
            begin
                // Must create 609/1024*Vdd
                Q = 30'b111110100000000000000000000000;
                prev_state = State0_609;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_305)
            begin
                // Must create 611/1024*Vdd
                Q = 30'b111000001100000000000000100000;
                prev_state = State0_611;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_307)
            begin
                // Must create 613/1024*Vdd
                Q = 30'b100000001100000000000000111000;
                prev_state = State0_613;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_307)
            begin
                // Must create 615/1024*Vdd
                Q = 30'b101000001100000000000000110000;
                prev_state = State0_615;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_309)
            begin
                // Must create 617/1024*Vdd
                Q = 30'b101100101000000000000000100000;
                prev_state = State0_617;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_309)
            begin
                // Must create 619/1024*Vdd
                Q = 30'b101100101100000000000000000000;
                prev_state = State0_619;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_311)
            begin
                // Must create 621/1024*Vdd
                Q = 30'b101100101100000000000000000000;
                prev_state = State0_621;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_311)
            begin
                // Must create 623/1024*Vdd
                Q = 30'b100000101100000000000100000001;
                prev_state = State0_623;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_313)
            begin
                // Must create 625/1024*Vdd
                Q = 30'b100010010000000000010000000000;
                prev_state = State0_625;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_313)
            begin
                // Must create 627/1024*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State0_627;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_315)
            begin
                // Must create 629/1024*Vdd
                Q = 30'b111100100000000001000000000000;
                prev_state = State0_629;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_315)
            begin
                // Must create 631/1024*Vdd
                Q = 30'b111100100000000000001000000000;
                prev_state = State0_631;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_317)
            begin
                // Must create 633/1024*Vdd
                Q = 30'b111011000000000001000000000000;
                prev_state = State0_633;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_317)
            begin
                // Must create 635/1024*Vdd
                Q = 30'b110011000000000001100000000000;
                prev_state = State0_635;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_319)
            begin
                // Must create 637/1024*Vdd
                Q = 30'b110011001000000100000000000000;
                prev_state = State0_637;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_319)
            begin
                // Must create 639/1024*Vdd
                Q = 30'b100000001000000000001100000000;
                prev_state = State0_639;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_321)
            begin
                // Must create 641/1024*Vdd
                Q = 30'b100000000000000000000100000000;
                prev_state = State0_641;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_321)
            begin
                // Must create 643/1024*Vdd
                Q = 30'b101000000000000000001100000000;
                prev_state = State0_643;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_323)
            begin
                // Must create 645/1024*Vdd
                Q = 30'b101000010000000010001100000000;
                prev_state = State0_645;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_323)
            begin
                // Must create 647/1024*Vdd
                Q = 30'b111000010000000000000100000001;
                prev_state = State0_647;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_325)
            begin
                // Must create 649/1024*Vdd
                Q = 30'b111000110000000000010000000000;
                prev_state = State0_649;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_325)
            begin
                // Must create 651/1024*Vdd
                Q = 30'b111000110000000100000000000000;
                prev_state = State0_651;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_327)
            begin
                // Must create 653/1024*Vdd
                Q = 30'b111000110000000100000000000000;
                prev_state = State0_653;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_327)
            begin
                // Must create 655/1024*Vdd
                Q = 30'b100001110000000100000000000001;
                prev_state = State0_655;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_329)
            begin
                // Must create 657/1024*Vdd
                Q = 30'b100000100000000100001000001100;
                prev_state = State0_657;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_329)
            begin
                // Must create 659/1024*Vdd
                Q = 30'b111000000000000100000000001100;
                prev_state = State0_659;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_331)
            begin
                // Must create 661/1024*Vdd
                Q = 30'b111000000000000100000000001100;
                prev_state = State0_661;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_331)
            begin
                // Must create 663/1024*Vdd
                Q = 30'b111000000000000100000000101000;
                prev_state = State0_663;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_333)
            begin
                // Must create 665/1024*Vdd
                Q = 30'b111010000000000100000000000100;
                prev_state = State0_665;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_333)
            begin
                // Must create 667/1024*Vdd
                Q = 30'b111010000000000100000000001000;
                prev_state = State0_667;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_335)
            begin
                // Must create 669/1024*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State0_669;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_335)
            begin
                // Must create 671/1024*Vdd
                Q = 30'b110000010000000000010000000011;
                prev_state = State0_671;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_337)
            begin
                // Must create 673/1024*Vdd
                Q = 30'b110010110000000000001000000000;
                prev_state = State0_673;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_337)
            begin
                // Must create 675/1024*Vdd
                Q = 30'b111101010000000000000000000000;
                prev_state = State0_675;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_339)
            begin
                // Must create 677/1024*Vdd
                Q = 30'b101101000000000000000000110000;
                prev_state = State0_677;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_339)
            begin
                // Must create 679/1024*Vdd
                Q = 30'b111101000000000000000000100000;
                prev_state = State0_679;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_341)
            begin
                // Must create 681/1024*Vdd
                Q = 30'b111111000000000000000000000000;
                prev_state = State0_681;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_341)
            begin
                // Must create 683/1024*Vdd
                Q = 30'b111110100000000000000000000000;
                prev_state = State0_683;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_343)
            begin
                // Must create 685/1024*Vdd
                Q = 30'b111110100000000000000000000000;
                prev_state = State0_685;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_343)
            begin
                // Must create 687/1024*Vdd
                Q = 30'b100110100000000000000010000001;
                prev_state = State0_687;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_345)
            begin
                // Must create 689/1024*Vdd
                Q = 30'b100011110000000000000000000001;
                prev_state = State0_689;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_345)
            begin
                // Must create 691/1024*Vdd
                Q = 30'b111010110000000000000000000000;
                prev_state = State0_691;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_347)
            begin
                // Must create 693/1024*Vdd
                Q = 30'b111010110000000000000000000000;
                prev_state = State0_693;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_347)
            begin
                // Must create 695/1024*Vdd
                Q = 30'b111010100000000001000000000000;
                prev_state = State0_695;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_349)
            begin
                // Must create 697/1024*Vdd
                Q = 30'b111000010000000000000001000001;
                prev_state = State0_697;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_349)
            begin
                // Must create 699/1024*Vdd
                Q = 30'b101000010000000000100011000000;
                prev_state = State0_699;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_351)
            begin
                // Must create 701/1024*Vdd
                Q = 30'b101000000000000000000011000000;
                prev_state = State0_701;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_351)
            begin
                // Must create 703/1024*Vdd
                Q = 30'b100000000000000000000001000000;
                prev_state = State0_703;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_353)
            begin
                // Must create 705/1024*Vdd
                Q = 30'b100000000000000000000001000000;
                prev_state = State0_705;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_353)
            begin
                // Must create 707/1024*Vdd
                Q = 30'b100000000000000001110101000000;
                prev_state = State0_707;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_355)
            begin
                // Must create 709/1024*Vdd
                Q = 30'b111000000000000000010100100000;
                prev_state = State0_709;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_355)
            begin
                // Must create 711/1024*Vdd
                Q = 30'b110010000000000000001000000000;
                prev_state = State0_711;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_357)
            begin
                // Must create 713/1024*Vdd
                Q = 30'b111000000000000001100010000000;
                prev_state = State0_713;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_357)
            begin
                // Must create 715/1024*Vdd
                Q = 30'b111000000000000001110000000000;
                prev_state = State0_715;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_359)
            begin
                // Must create 717/1024*Vdd
                Q = 30'b111000000000000001110000000000;
                prev_state = State0_717;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_359)
            begin
                // Must create 719/1024*Vdd
                Q = 30'b100000000000000101000110010000;
                prev_state = State0_719;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_361)
            begin
                // Must create 721/1024*Vdd
                Q = 30'b100100000000000100001010010000;
                prev_state = State0_721;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_361)
            begin
                // Must create 723/1024*Vdd
                Q = 30'b111100000000000100001000000000;
                prev_state = State0_723;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_363)
            begin
                // Must create 725/1024*Vdd
                Q = 30'b111110000000000001000000000000;
                prev_state = State0_725;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_363)
            begin
                // Must create 727/1024*Vdd
                Q = 30'b111000000000000001000000110000;
                prev_state = State0_727;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_365)
            begin
                // Must create 729/1024*Vdd
                Q = 30'b110100000000000100000011000000;
                prev_state = State0_729;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_365)
            begin
                // Must create 731/1024*Vdd
                Q = 30'b100100000000000100000011001000;
                prev_state = State0_731;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_367)
            begin
                // Must create 733/1024*Vdd
                Q = 30'b100100000000000010000011100000;
                prev_state = State0_733;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_367)
            begin
                // Must create 735/1024*Vdd
                Q = 30'b100000000000000000000000100000;
                prev_state = State0_735;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_369)
            begin
                // Must create 737/1024*Vdd
                Q = 30'b100000000000000000000000100000;
                prev_state = State0_737;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_369)
            begin
                // Must create 739/1024*Vdd
                Q = 30'b100000000000000100101010100000;
                prev_state = State0_739;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_371)
            begin
                // Must create 741/1024*Vdd
                Q = 30'b111000000000000000001010001000;
                prev_state = State0_741;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_371)
            begin
                // Must create 743/1024*Vdd
                Q = 30'b111000000000000000001011000000;
                prev_state = State0_743;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_373)
            begin
                // Must create 745/1024*Vdd
                Q = 30'b111010000000000000000011000000;
                prev_state = State0_745;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_373)
            begin
                // Must create 747/1024*Vdd
                Q = 30'b111000000000000000000011010000;
                prev_state = State0_747;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_375)
            begin
                // Must create 749/1024*Vdd
                Q = 30'b111000000000000000000011010000;
                prev_state = State0_749;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_375)
            begin
                // Must create 751/1024*Vdd
                Q = 30'b100010000000000100000010101000;
                prev_state = State0_751;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_377)
            begin
                // Must create 753/1024*Vdd
                Q = 30'b101000000000000000000011011000;
                prev_state = State0_753;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_377)
            begin
                // Must create 755/1024*Vdd
                Q = 30'b110000000000000001000011010000;
                prev_state = State0_755;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_379)
            begin
                // Must create 757/1024*Vdd
                Q = 30'b100000000000000001010011010000;
                prev_state = State0_757;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_379)
            begin
                // Must create 759/1024*Vdd
                Q = 30'b100000000000000001110011000000;
                prev_state = State0_759;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_381)
            begin
                // Must create 761/1024*Vdd
                Q = 30'b100000000000000101100010001000;
                prev_state = State0_761;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_381)
            begin
                // Must create 763/1024*Vdd
                Q = 30'b100000000000000101111000000000;
                prev_state = State0_763;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_383)
            begin
                // Must create 765/1024*Vdd
                Q = 30'b100000000000000111110000000000;
                prev_state = State0_765;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_383)
            begin
                // Must create 767/1024*Vdd
                Q = 30'b100000000000000000100000000000;
                prev_state = State0_767;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_385)
            begin
                // Must create 769/1024*Vdd
                Q = 30'b100000000000000000100000000000;
                prev_state = State0_769;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_385)
            begin
                // Must create 771/1024*Vdd
                Q = 30'b100100000000000001100000000000;
                prev_state = State0_771;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_387)
            begin
                // Must create 773/1024*Vdd
                Q = 30'b110000000000000000000000000000;
                prev_state = State0_773;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_387)
            begin
                // Must create 775/1024*Vdd
                Q = 30'b100000000000000000000000000010;
                prev_state = State0_775;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_389)
            begin
                // Must create 777/1024*Vdd
                Q = 30'b110100000000000000100000000110;
                prev_state = State0_777;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_389)
            begin
                // Must create 779/1024*Vdd
                Q = 30'b110100000000000110000000000100;
                prev_state = State0_779;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_391)
            begin
                // Must create 781/1024*Vdd
                Q = 30'b110100000000000110010000000000;
                prev_state = State0_781;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_391)
            begin
                // Must create 783/1024*Vdd
                Q = 30'b100000000000000110010000010010;
                prev_state = State0_783;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_393)
            begin
                // Must create 785/1024*Vdd
                Q = 30'b100000000000000100110000110000;
                prev_state = State0_785;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_393)
            begin
                // Must create 787/1024*Vdd
                Q = 30'b110100000000000100010000100000;
                prev_state = State0_787;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_395)
            begin
                // Must create 789/1024*Vdd
                Q = 30'b110100000000000100010000000100;
                prev_state = State0_789;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_395)
            begin
                // Must create 791/1024*Vdd
                Q = 30'b100000000000000000000000010000;
                prev_state = State0_791;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_397)
            begin
                // Must create 793/1024*Vdd
                Q = 30'b111100000000000100000000000100;
                prev_state = State0_793;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_397)
            begin
                // Must create 795/1024*Vdd
                Q = 30'b111100000000000100000000001000;
                prev_state = State0_795;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_399)
            begin
                // Must create 797/1024*Vdd
                Q = 30'b111100000000000000011000000000;
                prev_state = State0_797;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_399)
            begin
                // Must create 799/1024*Vdd
                Q = 30'b110000000000000001100110000000;
                prev_state = State0_799;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_401)
            begin
                // Must create 801/1024*Vdd
                Q = 30'b101000000000000000000000011000;
                prev_state = State0_801;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_401)
            begin
                // Must create 803/1024*Vdd
                Q = 30'b111100000000000101000000000000;
                prev_state = State0_803;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_403)
            begin
                // Must create 805/1024*Vdd
                Q = 30'b110100000000000001100000000100;
                prev_state = State0_805;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_403)
            begin
                // Must create 807/1024*Vdd
                Q = 30'b110100000000000001100000000010;
                prev_state = State0_807;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_405)
            begin
                // Must create 809/1024*Vdd
                Q = 30'b110100000000000001000000010100;
                prev_state = State0_809;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_405)
            begin
                // Must create 811/1024*Vdd
                Q = 30'b110100000000000001000000000110;
                prev_state = State0_811;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_407)
            begin
                // Must create 813/1024*Vdd
                Q = 30'b111000000000000001000000000110;
                prev_state = State0_813;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_407)
            begin
                // Must create 815/1024*Vdd
                Q = 30'b100000000000000001001000100110;
                prev_state = State0_815;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_409)
            begin
                // Must create 817/1024*Vdd
                Q = 30'b100000000000000101011000000100;
                prev_state = State0_817;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_409)
            begin
                // Must create 819/1024*Vdd
                Q = 30'b111000000000000101000000000100;
                prev_state = State0_819;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_411)
            begin
                // Must create 821/1024*Vdd
                Q = 30'b111000000000000101000000000010;
                prev_state = State0_821;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_411)
            begin
                // Must create 823/1024*Vdd
                Q = 30'b111000000000000000001010000010;
                prev_state = State0_823;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_413)
            begin
                // Must create 825/1024*Vdd
                Q = 30'b100000000000000000001000000000;
                prev_state = State0_825;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_413)
            begin
                // Must create 827/1024*Vdd
                Q = 30'b100000000000000000000100000000;
                prev_state = State0_827;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_415)
            begin
                // Must create 829/1024*Vdd
                Q = 30'b110000000000000000000011000000;
                prev_state = State0_829;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_415)
            begin
                // Must create 831/1024*Vdd
                Q = 30'b100000000000000000000001000000;
                prev_state = State0_831;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_417)
            begin
                // Must create 833/1024*Vdd
                Q = 30'b100000000000000000000001000000;
                prev_state = State0_833;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_417)
            begin
                // Must create 835/1024*Vdd
                Q = 30'b100000000000000000100101110000;
                prev_state = State0_835;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_419)
            begin
                // Must create 837/1024*Vdd
                Q = 30'b111000000000000000000000111000;
                prev_state = State0_837;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_419)
            begin
                // Must create 839/1024*Vdd
                Q = 30'b110000000000000001001000000000;
                prev_state = State0_839;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_421)
            begin
                // Must create 841/1024*Vdd
                Q = 30'b111000000000000000000110010000;
                prev_state = State0_841;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_421)
            begin
                // Must create 843/1024*Vdd
                Q = 30'b111000000000000000000100011000;
                prev_state = State0_843;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_423)
            begin
                // Must create 845/1024*Vdd
                Q = 30'b111000000000000000000100011000;
                prev_state = State0_845;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_423)
            begin
                // Must create 847/1024*Vdd
                Q = 30'b100000000000000010000110000110;
                prev_state = State0_847;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_425)
            begin
                // Must create 849/1024*Vdd
                Q = 30'b100000000000000000000000001000;
                prev_state = State0_849;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_425)
            begin
                // Must create 851/1024*Vdd
                Q = 30'b100000000000000101111000000000;
                prev_state = State0_851;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_427)
            begin
                // Must create 853/1024*Vdd
                Q = 30'b110000000000000100011000001000;
                prev_state = State0_853;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_427)
            begin
                // Must create 855/1024*Vdd
                Q = 30'b111000000000000100000000011000;
                prev_state = State0_855;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_429)
            begin
                // Must create 857/1024*Vdd
                Q = 30'b110000000000000010000001000011;
                prev_state = State0_857;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_429)
            begin
                // Must create 859/1024*Vdd
                Q = 30'b100000000000000101000001001100;
                prev_state = State0_859;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_431)
            begin
                // Must create 861/1024*Vdd
                Q = 30'b111000000000000000000011001000;
                prev_state = State0_861;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_431)
            begin
                // Must create 863/1024*Vdd
                Q = 30'b100000000000000000000000100000;
                prev_state = State0_863;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_433)
            begin
                // Must create 865/1024*Vdd
                Q = 30'b100000000000000000000000100000;
                prev_state = State0_865;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_433)
            begin
                // Must create 867/1024*Vdd
                Q = 30'b111000000000000100001001000000;
                prev_state = State0_867;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_435)
            begin
                // Must create 869/1024*Vdd
                Q = 30'b111000000000000101000010000000;
                prev_state = State0_869;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_435)
            begin
                // Must create 871/1024*Vdd
                Q = 30'b111000000000000101001000000000;
                prev_state = State0_871;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_437)
            begin
                // Must create 873/1024*Vdd
                Q = 30'b111000000000000101000000100000;
                prev_state = State0_873;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_437)
            begin
                // Must create 875/1024*Vdd
                Q = 30'b111000000000000101001000000000;
                prev_state = State0_875;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_439)
            begin
                // Must create 877/1024*Vdd
                Q = 30'b111000000000000101001000000000;
                prev_state = State0_877;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_439)
            begin
                // Must create 879/1024*Vdd
                Q = 30'b110000000000000000000100010000;
                prev_state = State0_879;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_441)
            begin
                // Must create 881/1024*Vdd
                Q = 30'b100000000000000000000000010000;
                prev_state = State0_881;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_441)
            begin
                // Must create 883/1024*Vdd
                Q = 30'b111000000000000000001011000000;
                prev_state = State0_883;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_443)
            begin
                // Must create 885/1024*Vdd
                Q = 30'b111000000000000000011010000000;
                prev_state = State0_885;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_443)
            begin
                // Must create 887/1024*Vdd
                Q = 30'b100000000000000001001100100100;
                prev_state = State0_887;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_445)
            begin
                // Must create 889/1024*Vdd
                Q = 30'b111000000000000000011000001000;
                prev_state = State0_889;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_445)
            begin
                // Must create 891/1024*Vdd
                Q = 30'b111000000000000001010010000000;
                prev_state = State0_891;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_447)
            begin
                // Must create 893/1024*Vdd
                Q = 30'b111000000000000001110000000000;
                prev_state = State0_893;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_447)
            begin
                // Must create 895/1024*Vdd
                Q = 30'b100000000000000000010000000000;
                prev_state = State0_895;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_449)
            begin
                // Must create 897/1024*Vdd
                Q = 30'b100000000000000000010000000000;
                prev_state = State0_897;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_449)
            begin
                // Must create 899/1024*Vdd
                Q = 30'b100000000000000110010000000110;
                prev_state = State0_899;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_451)
            begin
                // Must create 901/1024*Vdd
                Q = 30'b010000000000000110000000000111;
                prev_state = State0_901;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_451)
            begin
                // Must create 903/1024*Vdd
                Q = 30'b010000000000000111000000000110;
                prev_state = State0_903;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_453)
            begin
                // Must create 905/1024*Vdd
                Q = 30'b110000000000000101101000000000;
                prev_state = State0_905;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_453)
            begin
                // Must create 907/1024*Vdd
                Q = 30'b010000000000000101101010000000;
                prev_state = State0_907;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_455)
            begin
                // Must create 909/1024*Vdd
                Q = 30'b010000000000000101101001000000;
                prev_state = State0_909;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_455)
            begin
                // Must create 911/1024*Vdd
                Q = 30'b010000000000000000000001000000;
                prev_state = State0_911;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_457)
            begin
                // Must create 913/1024*Vdd
                Q = 30'b100000000000000001100000011100;
                prev_state = State0_913;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_457)
            begin
                // Must create 915/1024*Vdd
                Q = 30'b110000000000000101001100000000;
                prev_state = State0_915;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_459)
            begin
                // Must create 917/1024*Vdd
                Q = 30'b110000000000000101001001000000;
                prev_state = State0_917;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_459)
            begin
                // Must create 919/1024*Vdd
                Q = 30'b110000000000000100000011010000;
                prev_state = State0_919;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_461)
            begin
                // Must create 921/1024*Vdd
                Q = 30'b100000000000000000010001111000;
                prev_state = State0_921;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_461)
            begin
                // Must create 923/1024*Vdd
                Q = 30'b110000000000000100000001000110;
                prev_state = State0_923;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_463)
            begin
                // Must create 925/1024*Vdd
                Q = 30'b110000000000000000100001100100;
                prev_state = State0_925;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_463)
            begin
                // Must create 927/1024*Vdd
                Q = 30'b100000000000000000000000001000;
                prev_state = State0_927;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_465)
            begin
                // Must create 929/1024*Vdd
                Q = 30'b100000000000000000000000001000;
                prev_state = State0_929;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_465)
            begin
                // Must create 931/1024*Vdd
                Q = 30'b100000000000000001011100000100;
                prev_state = State0_931;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_467)
            begin
                // Must create 933/1024*Vdd
                Q = 30'b110000000000000100000100000110;
                prev_state = State0_933;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_467)
            begin
                // Must create 935/1024*Vdd
                Q = 30'b110000000000000000000000110000;
                prev_state = State0_935;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_469)
            begin
                // Must create 937/1024*Vdd
                Q = 30'b100000000000000000000000010000;
                prev_state = State0_937;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_469)
            begin
                // Must create 939/1024*Vdd
                Q = 30'b110000000000000100001001000100;
                prev_state = State0_939;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_471)
            begin
                // Must create 941/1024*Vdd
                Q = 30'b110000000000000100001001100000;
                prev_state = State0_941;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_471)
            begin
                // Must create 943/1024*Vdd
                Q = 30'b100000000000000000001011110000;
                prev_state = State0_943;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_473)
            begin
                // Must create 945/1024*Vdd
                Q = 30'b100000000000000000000000000100;
                prev_state = State0_945;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_473)
            begin
                // Must create 947/1024*Vdd
                Q = 30'b110000000000000100001001100000;
                prev_state = State0_947;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_475)
            begin
                // Must create 949/1024*Vdd
                Q = 30'b110000000000000100001100100000;
                prev_state = State0_949;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_475)
            begin
                // Must create 951/1024*Vdd
                Q = 30'b110000000000000100000010100010;
                prev_state = State0_951;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_477)
            begin
                // Must create 953/1024*Vdd
                Q = 30'b110000000000000000000001000010;
                prev_state = State0_953;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_477)
            begin
                // Must create 955/1024*Vdd
                Q = 30'b110000000000000100000000001101;
                prev_state = State0_955;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_479)
            begin
                // Must create 957/1024*Vdd
                Q = 30'b100000000000000000000010111100;
                prev_state = State0_957;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_479)
            begin
                // Must create 959/1024*Vdd
                Q = 30'b100000000000000000000010000000;
                prev_state = State0_959;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_481)
            begin
                // Must create 961/1024*Vdd
                Q = 30'b100000000000000000000010000000;
                prev_state = State0_961;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_481)
            begin
                // Must create 963/1024*Vdd
                Q = 30'b100000000000000000010010101100;
                prev_state = State0_963;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_483)
            begin
                // Must create 965/1024*Vdd
                Q = 30'b110000000000000001000000001110;
                prev_state = State0_965;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_483)
            begin
                // Must create 967/1024*Vdd
                Q = 30'b110000000000000000000001010000;
                prev_state = State0_967;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_485)
            begin
                // Must create 969/1024*Vdd
                Q = 30'b110000000000000001000010011000;
                prev_state = State0_969;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_485)
            begin
                // Must create 971/1024*Vdd
                Q = 30'b110000000000000001001100001000;
                prev_state = State0_971;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_487)
            begin
                // Must create 973/1024*Vdd
                Q = 30'b110000000000000001001001001000;
                prev_state = State0_973;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_487)
            begin
                // Must create 975/1024*Vdd
                Q = 30'b100000000000000000000000000010;
                prev_state = State0_975;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_489)
            begin
                // Must create 977/1024*Vdd
                Q = 30'b010000000000000000000000000010;
                prev_state = State0_977;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_489)
            begin
                // Must create 979/1024*Vdd
                Q = 30'b010000000000000001001100011000;
                prev_state = State0_979;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_491)
            begin
                // Must create 981/1024*Vdd
                Q = 30'b010000000000000001001100010010;
                prev_state = State0_981;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_491)
            begin
                // Must create 983/1024*Vdd
                Q = 30'b010000000000000001001001000011;
                prev_state = State0_983;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_493)
            begin
                // Must create 985/1024*Vdd
                Q = 30'b010000000000000001000001100011;
                prev_state = State0_985;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_493)
            begin
                // Must create 987/1024*Vdd
                Q = 30'b010000000000000001000001111000;
                prev_state = State0_987;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_495)
            begin
                // Must create 989/1024*Vdd
                Q = 30'b010000000000000001000001100000;
                prev_state = State0_989;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_495)
            begin
                // Must create 991/1024*Vdd
                Q = 30'b010000000000000000000000100000;
                prev_state = State0_991;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_497)
            begin
                // Must create 993/1024*Vdd
                Q = 30'b100000000000000000000000100000;
                prev_state = State0_993;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_497)
            begin
                // Must create 995/1024*Vdd
                Q = 30'b110000000000000000001101010000;
                prev_state = State0_995;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_499)
            begin
                // Must create 997/1024*Vdd
                Q = 30'b010000000000000000001101000000;
                prev_state = State0_997;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_499)
            begin
                // Must create 999/1024*Vdd
                Q = 30'b010000000000000000000110100110;
                prev_state = State0_999;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_501)
            begin
                // Must create 1001/1024*Vdd
                Q = 30'b010000000000000000001111010000;
                prev_state = State0_1001;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_501)
            begin
                // Must create 1003/1024*Vdd
                Q = 30'b010000000000000000001110010100;
                prev_state = State0_1003;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_503)
            begin
                // Must create 1005/1024*Vdd
                Q = 30'b010000000000000000000000000100;
                prev_state = State0_1005;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_503)
            begin
                // Must create 1007/1024*Vdd
                Q = 30'b010000000000000000001001000001;
                prev_state = State0_1007;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_505)
            begin
                // Must create 1009/1024*Vdd
                Q = 30'b010000000000000000001000100001;
                prev_state = State0_1009;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_505)
            begin
                // Must create 1011/1024*Vdd
                Q = 30'b010000000000000000000000000100;
                prev_state = State0_1011;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_507)
            begin
                // Must create 1013/1024*Vdd
                Q = 30'b010000000000000000001000001100;
                prev_state = State0_1013;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_507)
            begin
                // Must create 1015/1024*Vdd
                Q = 30'b010000000000000000001000011101;
                prev_state = State0_1015;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_509)
            begin
                // Must create 1017/1024*Vdd
                Q = 30'b010000000000000000000000001000;
                prev_state = State0_1017;
            end
        else if (comp_reg == 1'b1 && prev_state_reg == State1_509)
            begin
                // Must create 1019/1024*Vdd
                Q = 30'b010000000000000000000000011001;
                prev_state = State0_1019;
            end
        else if (comp_reg == 1'b0 && prev_state_reg == State1_511)
            begin
                // Must create 1021/1024*Vdd
                Q = 30'b010000000000000000000000001011;
                prev_state = State0_1021;
            end
        else
            begin
                // Must create 1023/1024*Vdd
                Q = 30'b010000000000000000000000000001;
                prev_state = State0_1023;
            end
    end
  endcase
  end
end
endmodule
